module dff(input clk, output q, input d);
endmodule
