// Author        : Matteo Lupi  <matteo.lupi@cern.ch>
//-----------------------------------------------------------------------------
// Description :
// This module is designed to target the import construct.
// The imported values are used in always_comb_import.sv.
// The purpose of the module is purely of testing.
//-----------------------------------------------------------------------------
// Date        Author  Note
// 2021.07.29  mlupi   Created
//-----------------------------------------------------------------------------

package my_package_pkg;
  parameter ZERO        = 1'b0;
  parameter TRUE        = 1'b1;
  parameter LSB_CNT_MAX = 3564;
endpackage
