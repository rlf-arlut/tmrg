module m4(i,o);
input i;
output o;
m1 instM1(.i(i),.o(o));
m3 instM3(.i(i),.o(o));
endmodule

