module a();
endmodule

module b();
    a a_inst ();
endmodule
