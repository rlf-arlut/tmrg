module notxor;
 reg x1;
 reg x2;
 wire x3=x1 ~^ x2;
endmodule
