module a;
    reg x = 5;
endmodule
