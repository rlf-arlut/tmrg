module for;
integer i;
reg x,y;

  

generate


for (i = 0; i < 16; i = i +1) begin
   assign	  x=1;
   integer s;

for (j = 0; i < 16; i = i +1) begin
   assign	  x=1;
end
end


endgenerate

endmodule
