module m2(i,o);
input i;
output o;
m1 instM1(.i(i),.o(o));
endmodule
