module c;
    parameter N=1;
    reg value = N;
endmodule
