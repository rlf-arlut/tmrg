module signed_literal;
    wire [3:0]a;
    wire [3:0]b;
    assign a = 4'sb0100;
    assign b = 4'b0100;
endmodule
