module test;
// tmrg default triplicate
// tmrg do_not_triplicate signal
reg    [13:0] signal [0:CLUST-1];
wire   [13:0] signal2;
assign signal2=signal;
endmodule

