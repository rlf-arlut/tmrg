module test;
/*
fds
fsd
fds
fds
*/
wire i;
// tmrg default
endmodule
