module test;
 reg y;
initial 
  begin: x
     y=1'b1;
  end
endmodule
