module test;
  function automatic mux;
    input a, b, c, d;
  endfunction
endmodule

