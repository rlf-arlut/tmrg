module comb01 (in,out);
  input in;
  output out;
  wire combFun;
  assign combLogic = ~in1;
  assign out = combLogic;
endmodule
