module m1(i,o);
input i;
output o;
endmodule
