module AN2HVTD0 (A1, A2, Z);
   input A1, A2;
   output Z;
endmodule
module AN2HVTD1 (A1, A2, Z);
   input A1, A2;
   output Z;
endmodule
module AN2HVTD2 (A1, A2, Z);
   input A1, A2;
   output Z;
endmodule
module AN2HVTD4 (A1, A2, Z);
   input A1, A2;
   output Z;
endmodule
module AN2HVTD8 (A1, A2, Z);
   input A1, A2;
   output Z;
endmodule
module AN2XHVTD1 (A1, A2, Z);
   input A1, A2;
   output Z;
endmodule
module AN3HVTD0 (A1, A2, A3, Z);
   input A1, A2, A3;
   output Z;
endmodule
module AN3HVTD1 (A1, A2, A3, Z);
   input A1, A2, A3;
   output Z;
endmodule
module AN3HVTD2 (A1, A2, A3, Z);
   input A1, A2, A3;
   output Z;
endmodule
module AN3HVTD4 (A1, A2, A3, Z);
   input A1, A2, A3;
   output Z;
endmodule
module AN3HVTD8 (A1, A2, A3, Z);
   input A1, A2, A3;
   output Z;
endmodule
module AN3XHVTD1 (A1, A2, A3, Z);
   input A1, A2, A3;
   output Z;
endmodule
module AN4HVTD0 (A1, A2, A3, A4, Z);
   input A1, A2, A3, A4;
   output Z;
endmodule
module AN4HVTD1 (A1, A2, A3, A4, Z);
   input A1, A2, A3, A4;
   output Z;
endmodule
module AN4HVTD2 (A1, A2, A3, A4, Z);
   input A1, A2, A3, A4;
   output Z;
endmodule
module AN4HVTD4 (A1, A2, A3, A4, Z);
   input A1, A2, A3, A4;
   output Z;
endmodule
module AN4HVTD8 (A1, A2, A3, A4, Z);
   input A1, A2, A3, A4;
   output Z;
endmodule
module AN4XHVTD1 (A1, A2, A3, A4, Z);
   input A1, A2, A3, A4;
   output Z;
endmodule
module ANTENNAHVT (I);
  input I;
endmodule
module AO211HVTD0 (A1, A2, B, C, Z);
   input A1, A2, B, C;
   output Z;
endmodule
module AO211HVTD1 (A1, A2, B, C, Z);
   input A1, A2, B, C;
   output Z;
endmodule
module AO211HVTD2 (A1, A2, B, C, Z);
   input A1, A2, B, C;
   output Z;
endmodule
module AO211HVTD4 (A1, A2, B, C, Z);
   input A1, A2, B, C;
   output Z;
endmodule
module AO21HVTD0 (A1, A2, B, Z);
   input A1, A2, B;
   output Z;
endmodule
module AO21HVTD1 (A1, A2, B, Z);
   input A1, A2, B;
   output Z;
endmodule
module AO21HVTD2 (A1, A2, B, Z);
   input A1, A2, B;
   output Z;
endmodule
module AO21HVTD4 (A1, A2, B, Z);
   input A1, A2, B;
   output Z;
endmodule
module AO221HVTD0 (A1, A2, B1, B2, C, Z);
   input A1, A2, B1, B2, C;
   output Z;
endmodule
module AO221HVTD1 (A1, A2, B1, B2, C, Z);
   input A1, A2, B1, B2, C;
   output Z;
endmodule
module AO221HVTD2 (A1, A2, B1, B2, C, Z);
   input A1, A2, B1, B2, C;
   output Z;
endmodule
module AO221HVTD4 (A1, A2, B1, B2, C, Z);
   input A1, A2, B1, B2, C;
   output Z;
endmodule
module AO222HVTD0 (A1, A2, B1, B2, C1, C2, Z);
   input A1, A2, B1, B2, C1, C2;
   output Z;
endmodule
module AO222HVTD1 (A1, A2, B1, B2, C1, C2, Z);
   input A1, A2, B1, B2, C1, C2;
   output Z;
endmodule
module AO222HVTD2 (A1, A2, B1, B2, C1, C2, Z);
   input A1, A2, B1, B2, C1, C2;
   output Z;
endmodule
module AO222HVTD4 (A1, A2, B1, B2, C1, C2, Z);
   input A1, A2, B1, B2, C1, C2;
   output Z;
endmodule
module AO22HVTD0 (A1, A2, B1, B2, Z);
   input A1, A2, B1, B2;
   output Z;
endmodule
module AO22HVTD1 (A1, A2, B1, B2, Z);
   input A1, A2, B1, B2;
   output Z;
endmodule
module AO22HVTD2 (A1, A2, B1, B2, Z);
   input A1, A2, B1, B2;
   output Z;
endmodule
module AO22HVTD4 (A1, A2, B1, B2, Z);
   input A1, A2, B1, B2;
   output Z;
endmodule
module AO31HVTD0 (A1, A2, A3, B, Z);
   input A1, A2, A3, B;
   output Z;
endmodule
module AO31HVTD1 (A1, A2, A3, B, Z);
   input A1, A2, A3, B;
   output Z;
endmodule
module AO31HVTD2 (A1, A2, A3, B, Z);
   input A1, A2, A3, B;
   output Z;
endmodule
module AO31HVTD4 (A1, A2, A3, B, Z);
   input A1, A2, A3, B;
   output Z;
endmodule
module AO32HVTD0 (A1, A2, A3, B1, B2, Z);
   input A1, A2, A3, B1, B2;
   output Z;
endmodule
module AO32HVTD1 (A1, A2, A3, B1, B2, Z);
   input A1, A2, A3, B1, B2;
   output Z;
endmodule
module AO32HVTD2 (A1, A2, A3, B1, B2, Z);
   input A1, A2, A3, B1, B2;
   output Z;
endmodule
module AO32HVTD4 (A1, A2, A3, B1, B2, Z);
   input A1, A2, A3, B1, B2;
   output Z;
endmodule
module AO33HVTD0 (A1, A2, A3, B1, B2, B3, Z);
   input A1, A2, A3, B1, B2, B3;
   output Z;
endmodule
module AO33HVTD1 (A1, A2, A3, B1, B2, B3, Z);
   input A1, A2, A3, B1, B2, B3;
   output Z;
endmodule
module AO33HVTD2 (A1, A2, A3, B1, B2, B3, Z);
   input A1, A2, A3, B1, B2, B3;
   output Z;
endmodule
module AO33HVTD4 (A1, A2, A3, B1, B2, B3, Z);
   input A1, A2, A3, B1, B2, B3;
   output Z;
endmodule
module AOI211HVTD0 (A1, A2, B, C, ZN);
   input A1, A2, B, C;
   output ZN;
endmodule
module AOI211HVTD1 (A1, A2, B, C, ZN);
   input A1, A2, B, C;
   output ZN;
endmodule
module AOI211HVTD2 (A1, A2, B, C, ZN);
   input A1, A2, B, C;
   output ZN;
endmodule
module AOI211HVTD4 (A1, A2, B, C, ZN);
   input A1, A2, B, C;
   output ZN;
endmodule
module AOI211XHVTD0 (A1, A2, B, C, ZN);
   input A1, A2, B, C;
   output ZN;
endmodule
module AOI211XHVTD1 (A1, A2, B, C, ZN);
   input A1, A2, B, C;
   output ZN;
endmodule
module AOI211XHVTD2 (A1, A2, B, C, ZN);
   input A1, A2, B, C;
   output ZN;
endmodule
module AOI211XHVTD4 (A1, A2, B, C, ZN);
   input A1, A2, B, C;
   output ZN;
endmodule
module AOI21HVTD0 (A1, A2, B, ZN);
   input A1, A2, B;
   output ZN;
endmodule
module AOI21HVTD1 (A1, A2, B, ZN);
   input A1, A2, B;
   output ZN;
endmodule
module AOI21HVTD2 (A1, A2, B, ZN);
   input A1, A2, B;
   output ZN;
endmodule
module AOI21HVTD4 (A1, A2, B, ZN);
   input A1, A2, B;
   output ZN;
endmodule
module AOI221HVTD0 (A1, A2, B1, B2, C, ZN);
   input A1, A2, B1, B2, C;
   output ZN;
endmodule
module AOI221HVTD1 (A1, A2, B1, B2, C, ZN);
   input A1, A2, B1, B2, C;
   output ZN;
endmodule
module AOI221HVTD2 (A1, A2, B1, B2, C, ZN);
   input A1, A2, B1, B2, C;
   output ZN;
endmodule
module AOI221HVTD4 (A1, A2, B1, B2, C, ZN);
   input A1, A2, B1, B2, C;
   output ZN;
endmodule
module AOI221XHVTD4 (A1, A2, B1, B2, C, ZN);
   input A1, A2, B1, B2, C;
   output ZN;
endmodule
module AOI222HVTD0 (A1, A2, B1, B2, C1, C2, ZN);
   input A1, A2, B1, B2, C1, C2;
   output ZN;
endmodule
module AOI222HVTD1 (A1, A2, B1, B2, C1, C2, ZN);
   input A1, A2, B1, B2, C1, C2;
   output ZN;
endmodule
module AOI222HVTD2 (A1, A2, B1, B2, C1, C2, ZN);
   input A1, A2, B1, B2, C1, C2;
   output ZN;
endmodule
module AOI222HVTD4 (A1, A2, B1, B2, C1, C2, ZN);
   input A1, A2, B1, B2, C1, C2;
   output ZN;
endmodule
module AOI222XHVTD4 (A1, A2, B1, B2, C1, C2, ZN);
   input A1, A2, B1, B2, C1, C2;
   output ZN;
endmodule
module AOI22HVTD0 (A1, A2, B1, B2, ZN);
   input A1, A2, B1, B2;
   output ZN;
endmodule
module AOI22HVTD1 (A1, A2, B1, B2, ZN);
   input A1, A2, B1, B2;
   output ZN;
endmodule
module AOI22HVTD2 (A1, A2, B1, B2, ZN);
   input A1, A2, B1, B2;
   output ZN;
endmodule
module AOI22HVTD4 (A1, A2, B1, B2, ZN);
   input A1, A2, B1, B2;
   output ZN;
endmodule
module AOI31HVTD0 (A1, A2, A3, B, ZN);
   input A1, A2, A3, B;
   output ZN;
endmodule
module AOI31HVTD1 (A1, A2, A3, B, ZN);
   input A1, A2, A3, B;
   output ZN;
endmodule
module AOI31HVTD2 (A1, A2, A3, B, ZN);
   input A1, A2, A3, B;
   output ZN;
endmodule
module AOI31HVTD4 (A1, A2, A3, B, ZN);
   input A1, A2, A3, B;
   output ZN;
endmodule
module AOI32HVTD0 (A1, A2, A3, B1, B2, ZN);
   input A1, A2, A3, B1, B2;
   output ZN;
endmodule
module AOI32HVTD1 (A1, A2, A3, B1, B2, ZN);
   input A1, A2, A3, B1, B2;
   output ZN;
endmodule
module AOI32HVTD2 (A1, A2, A3, B1, B2, ZN);
   input A1, A2, A3, B1, B2;
   output ZN;
endmodule
module AOI32HVTD4 (A1, A2, A3, B1, B2, ZN);
   input A1, A2, A3, B1, B2;
   output ZN;
endmodule
module AOI32XHVTD4 (A1, A2, A3, B1, B2, ZN);
   input A1, A2, A3, B1, B2;
   output ZN;
endmodule
module AOI33HVTD0 (A1, A2, A3, B1, B2, B3, ZN);
   input A1, A2, A3, B1, B2, B3;
   output ZN;
endmodule
module AOI33HVTD1 (A1, A2, A3, B1, B2, B3, ZN);
   input A1, A2, A3, B1, B2, B3;
   output ZN;
endmodule
module AOI33HVTD2 (A1, A2, A3, B1, B2, B3, ZN);
   input A1, A2, A3, B1, B2, B3;
   output ZN;
endmodule
module AOI33HVTD4 (A1, A2, A3, B1, B2, B3, ZN);
   input A1, A2, A3, B1, B2, B3;
   output ZN;
endmodule
module AOI33XHVTD4 (A1, A2, A3, B1, B2, B3, ZN);
   input A1, A2, A3, B1, B2, B3;
   output ZN;
endmodule
module BENCHVTD1 (M0, M1, M2, X2, A, S);
   input M0, M1, M2;
   output X2;
   output A ;
   output S ;
endmodule
module BENCHVTD2 (M0, M1, M2, X2, A, S);
   input M0, M1, M2;
   output X2;
   output A ;
   output S ;
endmodule
module BENCHVTD4 (M0, M1, M2, X2, A, S);
   input M0, M1, M2;
   output X2;
   output A ;
   output S ;
endmodule
module BHDHVT (Z);
endmodule
module BMLHVTD1 (X2, A, S, M0, M1, PP);
   input X2, A, S, M0, M1;
   output PP;
endmodule
module BMLHVTD2 (X2, A, S, M0, M1, PP);
   input X2, A, S, M0, M1;
   output PP;
endmodule
module BMLHVTD4 (X2, A, S, M0, M1, PP);
   input X2, A, S, M0, M1;
   output PP;
endmodule
module BUFFHVTD0 (I, Z);
   input I;
   output Z;
endmodule
module BUFFHVTD1 (I, Z);
   input I;
   output Z;
endmodule
module BUFFHVTD12 (I, Z);
   input I;
   output Z;
endmodule
module BUFFHVTD16 (I, Z);
   input I;
   output Z;
endmodule
module BUFFHVTD2 (I, Z);
   input I;
   output Z;
endmodule
module BUFFHVTD20 (I, Z);
   input I;
   output Z;
endmodule
module BUFFHVTD24 (I, Z);
   input I;
   output Z;
endmodule
module BUFFHVTD3 (I, Z);
   input I;
   output Z;
endmodule
module BUFFHVTD4 (I, Z);
   input I;
   output Z;
endmodule
module BUFFHVTD6 (I, Z);
   input I;
   output Z;
endmodule
module BUFFHVTD8 (I, Z);
   input I;
   output Z;
endmodule
module BUFTHVTD0 (I, OE, Z);
   input I, OE;
   output Z;
endmodule
module BUFTHVTD1 (I, OE, Z);
   input I, OE;
   output Z;
endmodule
module BUFTHVTD12 (I, OE, Z);
   input I, OE;
   output Z;
endmodule
module BUFTHVTD16 (I, OE, Z);
   input I, OE;
   output Z;
endmodule
module BUFTHVTD2 (I, OE, Z);
   input I, OE;
   output Z;
endmodule
module BUFTHVTD20 (I, OE, Z);
   input I, OE;
   output Z;
endmodule
module BUFTHVTD24 (I, OE, Z);
   input I, OE;
   output Z;
endmodule
module BUFTHVTD3 (I, OE, Z);
   input I, OE;
   output Z;
endmodule
module BUFTHVTD4 (I, OE, Z);
   input I, OE;
   output Z;
endmodule
module BUFTHVTD6 (I, OE, Z);
   input I, OE;
   output Z;
endmodule
module BUFTHVTD8 (I, OE, Z);
   input I, OE;
   output Z;
endmodule
module CKAN2HVTD0 (A1, A2, Z);
   input A1, A2;
   output Z;
endmodule
module CKAN2HVTD1 (A1, A2, Z);
   input A1, A2;
   output Z;
endmodule
module CKAN2HVTD2 (A1, A2, Z);
   input A1, A2;
   output Z;
endmodule
module CKAN2HVTD4 (A1, A2, Z);
   input A1, A2;
   output Z;
endmodule
module CKAN2HVTD8 (A1, A2, Z);
   input A1, A2;
   output Z;
endmodule
module CKBHVTD0 (CLK, C);
   input CLK;
   output C;
endmodule
module CKBHVTD1 (CLK, C);
   input CLK;
   output C;
endmodule
module CKBHVTD12 (CLK, C);
   input CLK;
   output C;
endmodule
module CKBHVTD16 (CLK, C);
   input CLK;
   output C;
endmodule
module CKBHVTD2 (CLK, C);
   input CLK;
   output C;
endmodule
module CKBHVTD20 (CLK, C);
   input CLK;
   output C;
endmodule
module CKBHVTD24 (CLK, C);
   input CLK;
   output C;
endmodule
module CKBHVTD3 (CLK, C);
   input CLK;
   output C;
endmodule
module CKBHVTD4 (CLK, C);
   input CLK;
   output C;
endmodule
module CKBHVTD6 (CLK, C);
   input CLK;
   output C;
endmodule
module CKBHVTD8 (CLK, C);
   input CLK;
   output C;
endmodule
module CKBXHVTD0 (I, Z);
   input I;
   output Z;
endmodule
module CKBXHVTD1 (I, Z);
   input I;
   output Z;
endmodule
module CKBXHVTD12 (I, Z);
   input I;
   output Z;
endmodule
module CKBXHVTD16 (I, Z);
   input I;
   output Z;
endmodule
module CKBXHVTD2 (I, Z);
   input I;
   output Z;
endmodule
module CKBXHVTD20 (I, Z);
   input I;
   output Z;
endmodule
module CKBXHVTD24 (I, Z);
   input I;
   output Z;
endmodule
module CKBXHVTD3 (I, Z);
   input I;
   output Z;
endmodule
module CKBXHVTD4 (I, Z);
   input I;
   output Z;
endmodule
module CKBXHVTD6 (I, Z);
   input I;
   output Z;
endmodule
module CKBXHVTD8 (I, Z);
   input I;
   output Z;
endmodule
module CKLHQHVTD1 ( Q, TE, CPN, E );
    input TE, CPN, E;
    output Q;
endmodule
module CKLHQHVTD12 ( Q, TE, CPN, E );
    input TE, CPN, E;
    output Q;
endmodule
module CKLHQHVTD16 ( Q, TE, CPN, E );
    input TE, CPN, E;
    output Q;
endmodule
module CKLHQHVTD2 ( Q, TE, CPN, E );
    input TE, CPN, E;
    output Q;
endmodule
module CKLHQHVTD20 ( Q, TE, CPN, E );
    input TE, CPN, E;
    output Q;
endmodule
module CKLHQHVTD24 ( Q, TE, CPN, E );
    input TE, CPN, E;
    output Q;
endmodule
module CKLHQHVTD3 ( Q, TE, CPN, E );
    input TE, CPN, E;
    output Q;
endmodule
module CKLHQHVTD4 ( Q, TE, CPN, E );
    input TE, CPN, E;
    output Q;
endmodule
module CKLHQHVTD6 ( Q, TE, CPN, E );
    input TE, CPN, E;
    output Q;
endmodule
module CKLHQHVTD8 ( Q, TE, CPN, E );
    input TE, CPN, E;
    output Q;
endmodule
module CKLNQHVTD1 (TE, E, CP, Q);
    input TE, E, CP;
    output Q;
endmodule
module CKLNQHVTD12 (TE, E, CP, Q);
    input TE, E, CP;
    output Q;
endmodule
module CKLNQHVTD16 (TE, E, CP, Q);
    input TE, E, CP;
    output Q;
endmodule
module CKLNQHVTD2 (TE, E, CP, Q);
    input TE, E, CP;
    output Q;
endmodule
module CKLNQHVTD20 (TE, E, CP, Q);
    input TE, E, CP;
    output Q;
endmodule
module CKLNQHVTD24 (TE, E, CP, Q);
    input TE, E, CP;
    output Q;
endmodule
module CKLNQHVTD3 (TE, E, CP, Q);
    input TE, E, CP;
    output Q;
endmodule
module CKLNQHVTD4 (TE, E, CP, Q);
    input TE, E, CP;
    output Q;
endmodule
module CKLNQHVTD6 (TE, E, CP, Q);
    input TE, E, CP;
    output Q;
endmodule
module CKLNQHVTD8 (TE, E, CP, Q);
    input TE, E, CP;
    output Q;
endmodule
module CKMUX2HVTD0 (I0, I1, S, Z);
   input I0, I1, S;
   output Z;
endmodule
module CKMUX2HVTD1 (I0, I1, S, Z);
   input I0, I1, S;
   output Z;
endmodule
module CKMUX2HVTD2 (I0, I1, S, Z);
   input I0, I1, S;
   output Z;
endmodule
module CKMUX2HVTD4 (I0, I1, S, Z);
   input I0, I1, S;
   output Z;
endmodule
module CKND2HVTD0 (A1, A2, ZN);
   input A1, A2;
   output ZN;
endmodule
module CKND2HVTD1 (A1, A2, ZN);
   input A1, A2;
   output ZN;
endmodule
module CKND2HVTD2 (A1, A2, ZN);
   input A1, A2;
   output ZN;
endmodule
module CKND2HVTD3 (A1, A2, ZN);
   input A1, A2;
   output ZN;
endmodule
module CKND2HVTD4 (A1, A2, ZN);
   input A1, A2;
   output ZN;
endmodule
module CKND2HVTD8 (A1, A2, ZN);
   input A1, A2;
   output ZN;
endmodule
module CKNHVTD0 (CLK, CN);
   input CLK;
   output CN;
endmodule
module CKNHVTD1 (CLK, CN);
   input CLK;
   output CN;
endmodule
module CKNHVTD12 (CLK, CN);
   input CLK;
   output CN;
endmodule
module CKNHVTD16 (CLK, CN);
   input CLK;
   output CN;
endmodule
module CKNHVTD2 (CLK, CN);
   input CLK;
   output CN;
endmodule
module CKNHVTD20 (CLK, CN);
   input CLK;
   output CN;
endmodule
module CKNHVTD24 (CLK, CN);
   input CLK;
   output CN;
endmodule
module CKNHVTD3 (CLK, CN);
   input CLK;
   output CN;
endmodule
module CKNHVTD4 (CLK, CN);
   input CLK;
   output CN;
endmodule
module CKNHVTD6 (CLK, CN);
   input CLK;
   output CN;
endmodule
module CKNHVTD8 (CLK, CN);
   input CLK;
   output CN;
endmodule
module CKNXHVTD0 (I, ZN);
    input I;
    output ZN;
endmodule
module CKNXHVTD1 (I, ZN);
    input I;
    output ZN;
endmodule
module CKNXHVTD12 (I, ZN);
    input I;
    output ZN;
endmodule
module CKNXHVTD16 (I, ZN);
    input I;
    output ZN;
endmodule
module CKNXHVTD2 (I, ZN);
    input I;
    output ZN;
endmodule
module CKNXHVTD20 (I, ZN);
    input I;
    output ZN;
endmodule
module CKNXHVTD24 (I, ZN);
    input I;
    output ZN;
endmodule
module CKNXHVTD3 (I, ZN);
    input I;
    output ZN;
endmodule
module CKNXHVTD4 (I, ZN);
    input I;
    output ZN;
endmodule
module CKNXHVTD6 (I, ZN);
    input I;
    output ZN;
endmodule
module CKNXHVTD8 (I, ZN);
    input I;
    output ZN;
endmodule
module CKXOR2HVTD0 (A1, A2, Z);
   input A1, A2;
   output Z;
endmodule
module CKXOR2HVTD1 (A1, A2, Z);
   input A1, A2;
   output Z;
endmodule
module CKXOR2HVTD2 (A1, A2, Z);
   input A1, A2;
   output Z;
endmodule
module CKXOR2HVTD4 (A1, A2, Z);
   input A1, A2;
   output Z;
endmodule
module CMPE22HVTD1 (A, B, S, CO);
input A, B;
output S, CO;
endmodule
module CMPE22HVTD2 (A, B, S, CO);
input A, B;
output S, CO;
endmodule
module CMPE32HVTD1 (A, B, CI, S, CO);
input A, B, CI;
output S, CO;
endmodule
module CMPE32HVTD2 (A, B, CI, S, CO);
input A, B, CI;
output S, CO;
endmodule
module CMPE42HVTD1 (A, B, C, D, CIX, S, COX, CO);
   input A, B, C, D, CIX;
   output S;
   output COX ;
   output CO ;
endmodule
module CMPE42HVTD2 (A, B, C, D, CIX, S, COX, CO);
   input A, B, C, D, CIX;
   output S;
   output COX ;
   output CO ;
endmodule
module DCAPHVT;
endmodule
module DCAPHVT16;
endmodule
module DCAPHVT32;
endmodule
module DCAPHVT4;
endmodule
module DCAPHVT64;
endmodule
module DCAPHVT8;
endmodule
module DELHVT0 (I, Z);
   input I;
   output Z;
endmodule
module DELHVT005 (I, Z);
   input I;
   output Z;
endmodule
module DELHVT01 (I, Z);
   input I;
   output Z;
endmodule
module DELHVT015 (I, Z);
   input I;
   output Z;
endmodule
module DELHVT02 (I, Z);
   input I;
   output Z;
endmodule
module DELHVT1 (I, Z);
   input I;
   output Z;
endmodule
module DELHVT2 (I, Z);
   input I;
   output Z;
endmodule
module DELHVT3 (I, Z);
   input I;
   output Z;
endmodule
module DELHVT4 (I, Z);
   input I;
   output Z;
endmodule
module DFCNHVTD1 (D, CP, CDN, Q, QN);
    input D, CP, CDN;
    output Q, QN;
endmodule
module DFCNHVTD2 (D, CP, CDN, Q, QN);
    input D, CP, CDN;
    output Q, QN;
endmodule
module DFCNHVTD4 (D, CP, CDN, Q, QN);
    input D, CP, CDN;
    output Q, QN;
endmodule
module DFCNQHVTD1 (D, CP, CDN, Q);
    input D, CP, CDN;
    output Q;
endmodule
module DFCNQHVTD2 (D, CP, CDN, Q);
    input D, CP, CDN;
    output Q;
endmodule
module DFCNQHVTD4 (D, CP, CDN, Q);
    input D, CP, CDN;
    output Q;
endmodule
module DFCSNHVTD1 (D, CP, CDN, SDN, Q, QN);
    input D, CP, CDN, SDN;
    output Q, QN;
endmodule
module DFCSNHVTD2 (D, CP, CDN, SDN, Q, QN);
    input D, CP, CDN, SDN;
    output Q, QN;
endmodule
module DFCSNHVTD4 (D, CP, CDN, SDN, Q, QN);
    input D, CP, CDN, SDN;
    output Q, QN;
endmodule
module DFCSNQHVTD1 (D, CP, CDN, SDN, Q);
    input D, CP, CDN, SDN;
    output Q;
endmodule
module DFCSNQHVTD2 (D, CP, CDN, SDN, Q);
    input D, CP, CDN, SDN;
    output Q;
endmodule
module DFCSNQHVTD4 (D, CP, CDN, SDN, Q);
    input D, CP, CDN, SDN;
    output Q;
endmodule
module DFHVTD1 (D, CP, Q, QN);
    input D, CP;
    output Q, QN;
endmodule
module DFHVTD2 (D, CP, Q, QN);
    input D, CP;
    output Q, QN;
endmodule
module DFHVTD4 (D, CP, Q, QN);
    input D, CP;
    output Q, QN;
endmodule
module DFKCNHVTD1 (D, CP, CN, Q, QN);
    input D, CP, CN;
    output Q, QN;
endmodule
module DFKCNHVTD2 (D, CP, CN, Q, QN);
    input D, CP, CN;
    output Q, QN;
endmodule
module DFKCNHVTD4 (D, CP, CN, Q, QN);
    input D, CP, CN;
    output Q, QN;
endmodule
module DFKCNQHVTD1 (D, CP, CN, Q);
    input D, CP, CN;
    output Q;
endmodule
module DFKCNQHVTD2 (D, CP, CN, Q);
    input D, CP, CN;
    output Q;
endmodule
module DFKCNQHVTD4 (D, CP, CN, Q);
    input D, CP, CN;
    output Q;
endmodule
module DFKCSNHVTD1 (D, CP, CN, SN, Q, QN);
    input D, CP, CN, SN;
    output Q, QN;
endmodule
module DFKCSNHVTD2 (D, CP, CN, SN, Q, QN);
    input D, CP, CN, SN;
    output Q, QN;
endmodule
module DFKCSNHVTD4 (D, CP, CN, SN, Q, QN);
    input D, CP, CN, SN;
    output Q, QN;
endmodule
module DFKSNHVTD1 (D, CP, SN, Q, QN);
    input D, CP, SN;
    output Q, QN;
endmodule
module DFKSNHVTD2 (D, CP, SN, Q, QN);
    input D, CP, SN;
    output Q, QN;
endmodule
module DFKSNHVTD4 (D, CP, SN, Q, QN);
    input D, CP, SN;
    output Q, QN;
endmodule
module DFNCNHVTD1 (D, CPN, CDN, Q, QN);
    input D, CPN, CDN;
    output Q, QN;
endmodule
module DFNCNHVTD2 (D, CPN, CDN, Q, QN);
    input D, CPN, CDN;
    output Q, QN;
endmodule
module DFNCNHVTD4 (D, CPN, CDN, Q, QN);
    input D, CPN, CDN;
    output Q, QN;
endmodule
module DFNCSNHVTD1 (D, CPN, CDN, SDN, Q, QN);
    input D, CPN, CDN, SDN;
    output Q, QN;
endmodule
module DFNCSNHVTD2 (D, CPN, CDN, SDN, Q, QN);
    input D, CPN, CDN, SDN;
    output Q, QN;
endmodule
module DFNCSNHVTD4 (D, CPN, CDN, SDN, Q, QN);
    input D, CPN, CDN, SDN;
    output Q, QN;
endmodule
module DFNHVTD1 (D, CPN, Q, QN);
    input D, CPN;
    output Q, QN;
endmodule
module DFNHVTD2 (D, CPN, Q, QN);
    input D, CPN;
    output Q, QN;
endmodule
module DFNHVTD4 (D, CPN, Q, QN);
    input D, CPN;
    output Q, QN;
endmodule
module DFNSNHVTD1 (D, CPN, SDN, Q, QN);
    input D, CPN, SDN;
    output Q, QN;
endmodule
module DFNSNHVTD2 (D, CPN, SDN, Q, QN);
    input D, CPN, SDN;
    output Q, QN;
endmodule
module DFNSNHVTD4 (D, CPN, SDN, Q, QN);
    input D, CPN, SDN;
    output Q, QN;
endmodule
module DFQHVTD1 (D, CP, Q);
    input D, CP;
    output Q;
endmodule
module DFQHVTD2 (D, CP, Q);
    input D, CP;
    output Q;
endmodule
module DFQHVTD4 (D, CP, Q);
    input D, CP;
    output Q;
endmodule
module DFSNHVTD1 (D, CP, SDN, Q, QN);
    input D, CP, SDN;
    output Q, QN;
endmodule
module DFSNHVTD2 (D, CP, SDN, Q, QN);
    input D, CP, SDN;
    output Q, QN;
endmodule
module DFSNHVTD4 (D, CP, SDN, Q, QN);
    input D, CP, SDN;
    output Q, QN;
endmodule
module DFSNQHVTD1 (D, CP, SDN, Q);
    input D, CP, SDN;
    output Q;
endmodule
module DFSNQHVTD2 (D, CP, SDN, Q);
    input D, CP, SDN;
    output Q;
endmodule
module DFSNQHVTD4 (D, CP, SDN, Q);
    input D, CP, SDN;
    output Q;
endmodule
module DFXHVTD1 (DA, DB, SA, CP, Q, QN);
    input DA, DB, SA, CP;
    output Q, QN;
endmodule
module DFXHVTD2 (DA, DB, SA, CP, Q, QN);
    input DA, DB, SA, CP;
    output Q, QN;
endmodule
module DFXHVTD4 (DA, DB, SA, CP, Q, QN);
    input DA, DB, SA, CP;
    output Q, QN;
endmodule
module DFXQHVTD1 (DA, DB, SA, CP, Q);
    input DA, DB, SA, CP;
    output Q;
endmodule
module DFXQHVTD2 (DA, DB, SA, CP, Q);
    input DA, DB, SA, CP;
    output Q;
endmodule
module DFXQHVTD4 (DA, DB, SA, CP, Q);
    input DA, DB, SA, CP;
    output Q;
endmodule
module EDFCNHVTD1 (D, E, CP, CDN, Q, QN);
    input D, E, CP, CDN;  
    output Q, QN;
endmodule
module EDFCNHVTD2 (D, E, CP, CDN, Q, QN);
    input D, E, CP, CDN;  
    output Q, QN;
endmodule
module EDFCNHVTD4 (D, E, CP, CDN, Q, QN);
    input D, E, CP, CDN;  
    output Q, QN;
endmodule
module EDFCNQHVTD1 (D, E, CP, CDN, Q);
    input D, E, CP, CDN;  
    output Q;
endmodule
module EDFCNQHVTD2 (D, E, CP, CDN, Q);
    input D, E, CP, CDN;  
    output Q;
endmodule
module EDFCNQHVTD4 (D, E, CP, CDN, Q);
    input D, E, CP, CDN;  
    output Q;
endmodule
module EDFHVTD1 (D, E, CP, Q, QN);
    input D, E, CP;  
    output Q, QN;
endmodule
module EDFHVTD2 (D, E, CP, Q, QN);
    input D, E, CP;  
    output Q, QN;
endmodule
module EDFHVTD4 (D, E, CP, Q, QN);
    input D, E, CP;  
    output Q, QN;
endmodule
module EDFKCNHVTD1 (D, E, CP, CN, Q, QN);
    input D, E, CP, CN;
    output Q, QN;
endmodule
module EDFKCNHVTD2 (D, E, CP, CN, Q, QN);
    input D, E, CP, CN;
    output Q, QN;
endmodule
module EDFKCNHVTD4 (D, E, CP, CN, Q, QN);
    input D, E, CP, CN;
    output Q, QN;
endmodule
module EDFKCNQHVTD1 (D, E, CP, CN, Q);
    input D, E, CP, CN;
    output Q;
endmodule
module EDFKCNQHVTD2 (D, E, CP, CN, Q);
    input D, E, CP, CN;
    output Q;
endmodule
module EDFKCNQHVTD4 (D, E, CP, CN, Q);
    input D, E, CP, CN;
    output Q;
endmodule
module EDFQHVTD1 (D, E, CP, Q);
    input D, E, CP;  
    output Q;
endmodule
module EDFQHVTD2 (D, E, CP, Q);
    input D, E, CP;  
    output Q;
endmodule
module EDFQHVTD4 (D, E, CP, Q);
    input D, E, CP;  
    output Q;
endmodule
module FA1HVTD0 (A, B, CI, S, CO);
  input		A, B, CI;
  output	S, CO;
endmodule
module FA1HVTD1 (A, B, CI, S, CO);
  input		A, B, CI;
  output	S, CO;
endmodule
module FA1HVTD2 (A, B, CI, S, CO);
  input		A, B, CI;
  output	S, CO;
endmodule
module FA1HVTD4 (A, B, CI, S, CO);
  input		A, B, CI;
  output	S, CO;
endmodule
module FCICINHVTD1 (A, B, CIN, CO);
input A, B, CIN;
output CO;
endmodule
module FCICINHVTD2 (A, B, CIN, CO);
input A, B, CIN;
output CO;
endmodule
module FCICONHVTD1 (A, B, CI, CON);
input A, B, CI;
output CON;
endmodule
module FCICONHVTD2 (A, B, CI, CON);
input A, B, CI;
output CON;
endmodule
module FCSICINHVTD1 (A, B, CIN0, CIN1, CS, S, CO0, CO1);
input A, B, CIN0, CIN1, CS;
output S, CO0, CO1;
endmodule
module FCSICINHVTD2 (A, B, CIN0, CIN1, CS, S, CO0, CO1);
input A, B, CIN0, CIN1, CS;
output S, CO0, CO1;
endmodule
module FCSICONHVTD1 (A, B, CI0, CI1, CS, S, CON0, CON1);
input A, B, CI0, CI1, CS;
output S, CON0, CON1;
endmodule
module FCSICONHVTD2 (A, B, CI0, CI1, CS, S, CON0, CON1);
input A, B, CI0, CI1, CS;
output S, CON0, CON1;
endmodule
module FICINHVTD1 (A, B, CIN, S, CO);
input A, B, CIN;
output S, CO;
endmodule
module FICINHVTD2 (A, B, CIN, S, CO);
input A, B, CIN;
output S, CO;
endmodule
module FICONHVTD1 (A, B, CI, S, CON);
input A, B, CI;
output S, CON;
endmodule
module FICONHVTD2 (A, B, CI, S, CON);
input A, B, CI;
output S, CON;
endmodule
module FIICONHVTD1 (A, B, C, S, CON0, CON1);
input A, B, C;
output S, CON0, CON1;
endmodule
module FIICONHVTD2 (A, B, C, S, CON0, CON1);
input A, B, C;
output S, CON0, CON1;
endmodule
module HA1HVTD0 (A, B, S, CO);
  input	 	A, B;
  output	S, CO;
endmodule
module HA1HVTD1 (A, B, S, CO);
  input	 	A, B;
  output	S, CO;
endmodule
module HA1HVTD2 (A, B, S, CO);
  input	 	A, B;
  output	S, CO;
endmodule
module HA1HVTD4 (A, B, S, CO);
  input	 	A, B;
  output	S, CO;
endmodule
module HCOSCINHVTD1 (A, CIN, CS, S, CO);
input A, CIN, CS;
output S, CO;
endmodule
module HCOSCINHVTD2 (A, CIN, CS, S, CO);
input A, CIN, CS;
output S, CO;
endmodule
module HCOSCONHVTD1 (A, CI, CS, S, CON);
input A, CI, CS;
output S, CON;
endmodule
module HCOSCONHVTD2 (A, CI, CS, S, CON);
input A, CI, CS;
output S, CON;
endmodule
module HICINHVTD1 (A, CIN, S, CO);
input A, CIN;
output S, CO;
endmodule
module HICINHVTD2 (A, CIN, S, CO);
input A, CIN;
output S, CO;
endmodule
module HICONHVTD1 (A, CI, S, CON);
input A, CI;
output S, CON;
endmodule
module HICONHVTD2 (A, CI, S, CON);
input A, CI;
output S, CON;
endmodule
module IAO21HVTD0 (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
endmodule
module IAO21HVTD1 (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
endmodule
module IAO21HVTD2 (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
endmodule
module IAO21HVTD4 (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
endmodule
module IAO22HVTD0 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
endmodule
module IAO22HVTD1 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
endmodule
module IAO22HVTD2 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
endmodule
module IAO22HVTD4 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
endmodule
module IIND4HVTD0 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
endmodule
module IIND4HVTD1 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
endmodule
module IIND4HVTD2 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
endmodule
module IIND4HVTD4 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
endmodule
module IINR4HVTD0 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
endmodule
module IINR4HVTD1 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
endmodule
module IINR4HVTD2 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
endmodule
module IINR4HVTD4 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
endmodule
module IND2HVTD0 (A1, B1, ZN);
    input A1, B1;
    output ZN;
endmodule
module IND2HVTD1 (A1, B1, ZN);
    input A1, B1;
    output ZN;
endmodule
module IND2HVTD2 (A1, B1, ZN);
    input A1, B1;
    output ZN;
endmodule
module IND2HVTD4 (A1, B1, ZN);
    input A1, B1;
    output ZN;
endmodule
module IND3HVTD0 (A1, B1, B2, ZN);
    input A1, B1, B2;
    output ZN;
endmodule
module IND3HVTD1 (A1, B1, B2, ZN);
    input A1, B1, B2;
    output ZN;
endmodule
module IND3HVTD2 (A1, B1, B2, ZN);
    input A1, B1, B2;
    output ZN;
endmodule
module IND3HVTD4 (A1, B1, B2, ZN);
    input A1, B1, B2;
    output ZN;
endmodule
module IND4HVTD0 (A1, B1, B2, B3, ZN);
    input A1, B1, B2, B3;
    output ZN;
endmodule
module IND4HVTD1 (A1, B1, B2, B3, ZN);
    input A1, B1, B2, B3;
    output ZN;
endmodule
module IND4HVTD2 (A1, B1, B2, B3, ZN);
    input A1, B1, B2, B3;
    output ZN;
endmodule
module IND4HVTD4 (A1, B1, B2, B3, ZN);
    input A1, B1, B2, B3;
    output ZN;
endmodule
module INR2HVTD0 (A1, B1, ZN);
    input A1, B1;
    output ZN;
endmodule
module INR2HVTD1 (A1, B1, ZN);
    input A1, B1;
    output ZN;
endmodule
module INR2HVTD2 (A1, B1, ZN);
    input A1, B1;
    output ZN;
endmodule
module INR2HVTD4 (A1, B1, ZN);
    input A1, B1;
    output ZN;
endmodule
module INR2XHVTD0 (A1, B1, ZN);
    input A1, B1;
    output ZN;
endmodule
module INR2XHVTD1 (A1, B1, ZN);
    input A1, B1;
    output ZN;
endmodule
module INR2XHVTD2 (A1, B1, ZN);
    input A1, B1;
    output ZN;
endmodule
module INR2XHVTD4 (A1, B1, ZN);
    input A1, B1;
    output ZN;
endmodule
module INR3HVTD0 (A1, B1, B2, ZN);
    input A1, B1, B2;
    output ZN;
endmodule
module INR3HVTD1 (A1, B1, B2, ZN);
    input A1, B1, B2;
    output ZN;
endmodule
module INR3HVTD2 (A1, B1, B2, ZN);
    input A1, B1, B2;
    output ZN;
endmodule
module INR3HVTD4 (A1, B1, B2, ZN);
    input A1, B1, B2;
    output ZN;
endmodule
module INR4HVTD0 (A1, B1, B2, B3, ZN);
    input A1, B1, B2, B3;
    output ZN;
endmodule
module INR4HVTD1 (A1, B1, B2, B3, ZN);
    input A1, B1, B2, B3;
    output ZN;
endmodule
module INR4HVTD2 (A1, B1, B2, B3, ZN);
    input A1, B1, B2, B3;
    output ZN;
endmodule
module INR4HVTD4 (A1, B1, B2, B3, ZN);
    input A1, B1, B2, B3;
    output ZN;
endmodule
module INVHVTD0 (I, ZN);
    input I;
    output ZN;
endmodule
module INVHVTD1 (I, ZN);
    input I;
    output ZN;
endmodule
module INVHVTD12 (I, ZN);
    input I;
    output ZN;
endmodule
module INVHVTD16 (I, ZN);
    input I;
    output ZN;
endmodule
module INVHVTD2 (I, ZN);
    input I;
    output ZN;
endmodule
module INVHVTD20 (I, ZN);
    input I;
    output ZN;
endmodule
module INVHVTD24 (I, ZN);
    input I;
    output ZN;
endmodule
module INVHVTD3 (I, ZN);
    input I;
    output ZN;
endmodule
module INVHVTD4 (I, ZN);
    input I;
    output ZN;
endmodule
module INVHVTD6 (I, ZN);
    input I;
    output ZN;
endmodule
module INVHVTD8 (I, ZN);
    input I;
    output ZN;
endmodule
module IOA21HVTD0 (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
endmodule
module IOA21HVTD1 (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
endmodule
module IOA21HVTD2 (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
endmodule
module IOA21HVTD4 (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
endmodule
module IOA22HVTD0 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
endmodule
module IOA22HVTD1 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
endmodule
module IOA22HVTD2 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
endmodule
module IOA22HVTD4 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
endmodule
module LHCNHVTD1 (D, E, CDN, Q, QN);
    input D, E, CDN;
    output Q, QN;
endmodule
module LHCNHVTD2 (D, E, CDN, Q, QN);
    input D, E, CDN;
    output Q, QN;
endmodule
module LHCNHVTD4 (D, E, CDN, Q, QN);
    input D, E, CDN;
    output Q, QN;
endmodule
module LHCNQHVTD1 (D, E, CDN, Q);
    input D, E, CDN;
    output Q;
endmodule
module LHCNQHVTD2 (D, E, CDN, Q);
    input D, E, CDN;
    output Q;
endmodule
module LHCNQHVTD4 (D, E, CDN, Q);
    input D, E, CDN;
    output Q;
endmodule
module LHCSNHVTD1 (D, E, CDN, SDN, Q, QN);
    input D, E, CDN, SDN;
    output Q, QN;
endmodule
module LHCSNHVTD2 (D, E, CDN, SDN, Q, QN);
    input D, E, CDN, SDN;
    output Q, QN;
endmodule
module LHCSNHVTD4 (D, E, CDN, SDN, Q, QN);
    input D, E, CDN, SDN;
    output Q, QN;
endmodule
module LHCSNQHVTD1 (D, E, CDN, SDN, Q);
    input D, E, CDN, SDN;
    output Q;
endmodule
module LHCSNQHVTD2 (D, E, CDN, SDN, Q);
    input D, E, CDN, SDN;
    output Q;
endmodule
module LHCSNQHVTD4 (D, E, CDN, SDN, Q);
    input D, E, CDN, SDN;
    output Q;
endmodule
module LHHVTD1 (D, E, Q, QN);
    input D, E;
    output Q, QN;
endmodule
module LHHVTD2 (D, E, Q, QN);
    input D, E;
    output Q, QN;
endmodule
module LHHVTD4 (D, E, Q, QN);
    input D, E;
    output Q, QN;
endmodule
module LHQHVTD1 (D, E, Q);
    input D, E;
    output Q;
endmodule
module LHQHVTD2 (D, E, Q);
    input D, E;
    output Q;
endmodule
module LHQHVTD4 (D, E, Q);
    input D, E;
    output Q;
endmodule
module LHSNHVTD1 (D, E, SDN, Q, QN);
    input D, E, SDN;
    output Q, QN;
endmodule
module LHSNHVTD2 (D, E, SDN, Q, QN);
    input D, E, SDN;
    output Q, QN;
endmodule
module LHSNHVTD4 (D, E, SDN, Q, QN);
    input D, E, SDN;
    output Q, QN;
endmodule
module LHSNQHVTD1 (D, E, SDN, Q);
    input D, E, SDN;
    output Q;
endmodule
module LHSNQHVTD2 (D, E, SDN, Q);
    input D, E, SDN;
    output Q;
endmodule
module LHSNQHVTD4 (D, E, SDN, Q);
    input D, E, SDN;
    output Q;
endmodule
module LNCNHVTD1 (D, EN, CDN, Q, QN);
    input D, EN, CDN;
    output Q, QN;
endmodule
module LNCNHVTD2 (D, EN, CDN, Q, QN);
    input D, EN, CDN;
    output Q, QN;
endmodule
module LNCNHVTD4 (D, EN, CDN, Q, QN);
    input D, EN, CDN;
    output Q, QN;
endmodule
module LNCNQHVTD1 (D, EN, CDN, Q);
    input D, EN, CDN;
    output Q;
endmodule
module LNCNQHVTD2 (D, EN, CDN, Q);
    input D, EN, CDN;
    output Q;
endmodule
module LNCNQHVTD4 (D, EN, CDN, Q);
    input D, EN, CDN;
    output Q;
endmodule
module LNCSNHVTD1 (D, EN, CDN, SDN, Q, QN);
   input D, EN, CDN, SDN;
   output Q, QN;
endmodule
module LNCSNHVTD2 (D, EN, CDN, SDN, Q, QN);
   input D, EN, CDN, SDN;
   output Q, QN;
endmodule
module LNCSNHVTD4 (D, EN, CDN, SDN, Q, QN);
   input D, EN, CDN, SDN;
   output Q, QN;
endmodule
module LNCSNQHVTD1 (D, EN, CDN, SDN, Q);
   input D, EN, CDN, SDN;
   output Q;
endmodule
module LNCSNQHVTD2 (D, EN, CDN, SDN, Q);
   input D, EN, CDN, SDN;
   output Q;
endmodule
module LNCSNQHVTD4 (D, EN, CDN, SDN, Q);
   input D, EN, CDN, SDN;
   output Q;
endmodule
module LNHVTD1 (D, EN, Q, QN);
    input D, EN;
    output Q, QN;
endmodule
module LNHVTD2 (D, EN, Q, QN);
    input D, EN;
    output Q, QN;
endmodule
module LNHVTD4 (D, EN, Q, QN);
    input D, EN;
    output Q, QN;
endmodule
module LNQHVTD1 (D, EN, Q);
    input D, EN;
    output Q;
endmodule
module LNQHVTD2 (D, EN, Q);
    input D, EN;
    output Q;
endmodule
module LNQHVTD4 (D, EN, Q);
    input D, EN;
    output Q;
endmodule
module LNSNHVTD1 (D, EN, SDN, Q, QN);
    input D, EN, SDN;
    output Q, QN;
endmodule
module LNSNHVTD2 (D, EN, SDN, Q, QN);
    input D, EN, SDN;
    output Q, QN;
endmodule
module LNSNHVTD4 (D, EN, SDN, Q, QN);
    input D, EN, SDN;
    output Q, QN;
endmodule
module LNSNQHVTD1 (D, EN, SDN, Q);
    input D, EN, SDN;
    output Q;
endmodule
module LNSNQHVTD2 (D, EN, SDN, Q);
    input D, EN, SDN;
    output Q;
endmodule
module LNSNQHVTD4 (D, EN, SDN, Q);
    input D, EN, SDN;
    output Q;
endmodule
module MAOI222HVTD0 (A, B, C, ZN);
    input A, B, C;
    output ZN;
endmodule
module MAOI222HVTD1 (A, B, C, ZN);
    input A, B, C;
    output ZN;
endmodule
module MAOI222HVTD2 (A, B, C, ZN);
    input A, B, C;
    output ZN;
endmodule
module MAOI222HVTD4 (A, B, C, ZN);
    input A, B, C;
    output ZN;
endmodule
module MAOI22HVTD0 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
endmodule
module MAOI22HVTD1 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
endmodule
module MAOI22HVTD2 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
endmodule
module MAOI22HVTD4 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
endmodule
module MOAI22HVTD0 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
endmodule
module MOAI22HVTD1 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
endmodule
module MOAI22HVTD2 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
endmodule
module MOAI22HVTD4 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
endmodule
module MUX2HVTD0 (I0, I1, S, Z);
  input		I0, I1, S;
  output	Z;
endmodule
module MUX2HVTD1 (I0, I1, S, Z);
  input		I0, I1, S;
  output	Z;
endmodule
module MUX2HVTD2 (I0, I1, S, Z);
  input		I0, I1, S;
  output	Z;
endmodule
module MUX2HVTD4 (I0, I1, S, Z);
  input		I0, I1, S;
  output	Z;
endmodule
module MUX2NHVTD0 (I0, I1, S, ZN);
  input		 I0, I1, S;
  output	 ZN;
endmodule
module MUX2NHVTD1 (I0, I1, S, ZN);
  input		 I0, I1, S;
  output	 ZN;
endmodule
module MUX2NHVTD2 (I0, I1, S, ZN);
  input		 I0, I1, S;
  output	 ZN;
endmodule
module MUX2NHVTD4 (I0, I1, S, ZN);
  input		 I0, I1, S;
  output	 ZN;
endmodule
module MUX3HVTD0 (I0, I1, I2, S0, S1, Z);
  input		I0, I1, I2, S0, S1;
  output	Z;
endmodule
module MUX3HVTD1 (I0, I1, I2, S0, S1, Z);
  input		I0, I1, I2, S0, S1;
  output	Z;
endmodule
module MUX3HVTD2 (I0, I1, I2, S0, S1, Z);
  input		I0, I1, I2, S0, S1;
  output	Z;
endmodule
module MUX3HVTD4 (I0, I1, I2, S0, S1, Z);
  input		I0, I1, I2, S0, S1;
  output	Z;
endmodule
module MUX3NHVTD0 (I0, I1, I2, S0, S1, ZN);
  input 	I0, I1, I2, S0, S1;
  output 	ZN;
endmodule
module MUX3NHVTD1 (I0, I1, I2, S0, S1, ZN);
  input 	I0, I1, I2, S0, S1;
  output 	ZN;
endmodule
module MUX3NHVTD2 (I0, I1, I2, S0, S1, ZN);
  input 	I0, I1, I2, S0, S1;
  output 	ZN;
endmodule
module MUX3NHVTD4 (I0, I1, I2, S0, S1, ZN);
  input 	I0, I1, I2, S0, S1;
  output 	ZN;
endmodule
module MUX4HVTD0 (I0, I1, I2, I3, S0, S1, Z);
  input		 I0, I1, I2, I3, S0, S1;
  output	 Z;
endmodule
module MUX4HVTD1 (I0, I1, I2, I3, S0, S1, Z);
  input		 I0, I1, I2, I3, S0, S1;
  output	 Z;
endmodule
module MUX4HVTD2 (I0, I1, I2, I3, S0, S1, Z);
  input		 I0, I1, I2, I3, S0, S1;
  output	 Z;
endmodule
module MUX4HVTD4 (I0, I1, I2, I3, S0, S1, Z);
  input		 I0, I1, I2, I3, S0, S1;
  output	 Z;
endmodule
module MUX4NHVTD0 (I0, I1, I2, I3, S0, S1, ZN);
  input		 I0, I1, I2, I3, S0, S1;
  output	 ZN;
endmodule
module MUX4NHVTD1 (I0, I1, I2, I3, S0, S1, ZN);
  input		 I0, I1, I2, I3, S0, S1;
  output	 ZN;
endmodule
module MUX4NHVTD2 (I0, I1, I2, I3, S0, S1, ZN);
  input		 I0, I1, I2, I3, S0, S1;
  output	 ZN;
endmodule
module MUX4NHVTD4 (I0, I1, I2, I3, S0, S1, ZN);
  input		 I0, I1, I2, I3, S0, S1;
  output	 ZN;
endmodule
module ND2HVTD0 (A1, A2, ZN);
    input A1, A2;
    output ZN;
endmodule
module ND2HVTD1 (A1, A2, ZN);
    input A1, A2;
    output ZN;
endmodule
module ND2HVTD2 (A1, A2, ZN);
    input A1, A2;
    output ZN;
endmodule
module ND2HVTD3 (A1, A2, ZN);
    input A1, A2;
    output ZN;
endmodule
module ND2HVTD4 (A1, A2, ZN);
    input A1, A2;
    output ZN;
endmodule
module ND2HVTD8 (A1, A2, ZN);
    input A1, A2;
    output ZN;
endmodule
module ND3HVTD0 (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
endmodule
module ND3HVTD1 (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
endmodule
module ND3HVTD2 (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
endmodule
module ND3HVTD3 (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
endmodule
module ND3HVTD4 (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
endmodule
module ND3HVTD8 (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
endmodule
module ND4HVTD0 (A1, A2, A3, A4, ZN);
    input A1, A2, A3, A4;
    output ZN;
endmodule
module ND4HVTD1 (A1, A2, A3, A4, ZN);
    input A1, A2, A3, A4;
    output ZN;
endmodule
module ND4HVTD2 (A1, A2, A3, A4, ZN);
    input A1, A2, A3, A4;
    output ZN;
endmodule
module ND4HVTD3 (A1, A2, A3, A4, ZN);
    input A1, A2, A3, A4;
    output ZN;
endmodule
module ND4HVTD4 (A1, A2, A3, A4, ZN);
    input A1, A2, A3, A4;
    output ZN;
endmodule
module ND4HVTD8 (A1, A2, A3, A4, ZN);
    input A1, A2, A3, A4;
    output ZN;
endmodule
module NR2HVTD0 (A1, A2, ZN);
    input A1, A2;
    output ZN;
endmodule
module NR2HVTD1 (A1, A2, ZN);
    input A1, A2;
    output ZN;
endmodule
module NR2HVTD2 (A1, A2, ZN);
    input A1, A2;
    output ZN;
endmodule
module NR2HVTD3 (A1, A2, ZN);
    input A1, A2;
    output ZN;
endmodule
module NR2HVTD4 (A1, A2, ZN);
    input A1, A2;
    output ZN;
endmodule
module NR2HVTD8 (A1, A2, ZN);
    input A1, A2;
    output ZN;
endmodule
module NR2XHVTD0 (A1, A2, ZN);
    input A1, A2;
    output ZN;
endmodule
module NR2XHVTD1 (A1, A2, ZN);
    input A1, A2;
    output ZN;
endmodule
module NR2XHVTD2 (A1, A2, ZN);
    input A1, A2;
    output ZN;
endmodule
module NR2XHVTD3 (A1, A2, ZN);
    input A1, A2;
    output ZN;
endmodule
module NR2XHVTD4 (A1, A2, ZN);
    input A1, A2;
    output ZN;
endmodule
module NR2XHVTD8 (A1, A2, ZN);
    input A1, A2;
    output ZN;
endmodule
module NR3HVTD0 (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
endmodule
module NR3HVTD1 (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
endmodule
module NR3HVTD2 (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
endmodule
module NR3HVTD3 (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
endmodule
module NR3HVTD4 (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
endmodule
module NR3HVTD8 (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
endmodule
module NR4HVTD0 (A1, A2, A3, A4, ZN);
    input A1, A2, A3, A4;
    output ZN;
endmodule
module NR4HVTD1 (A1, A2, A3, A4, ZN);
    input A1, A2, A3, A4;
    output ZN;
endmodule
module NR4HVTD2 (A1, A2, A3, A4, ZN);
    input A1, A2, A3, A4;
    output ZN;
endmodule
module NR4HVTD3 (A1, A2, A3, A4, ZN);
    input A1, A2, A3, A4;
    output ZN;
endmodule
module NR4HVTD4 (A1, A2, A3, A4, ZN);
    input A1, A2, A3, A4;
    output ZN;
endmodule
module NR4HVTD8 (A1, A2, A3, A4, ZN);
    input A1, A2, A3, A4;
    output ZN;
endmodule
module OA211HVTD0 (A1, A2, B, C, Z);
    input A1, A2, B, C;
    output Z;
endmodule
module OA211HVTD1 (A1, A2, B, C, Z);
    input A1, A2, B, C;
    output Z;
endmodule
module OA211HVTD2 (A1, A2, B, C, Z);
    input A1, A2, B, C;
    output Z;
endmodule
module OA211HVTD4 (A1, A2, B, C, Z);
    input A1, A2, B, C;
    output Z;
endmodule
module OA21HVTD0 (A1, A2, B, Z);
    input A1, A2, B;
    output Z;
endmodule
module OA21HVTD1 (A1, A2, B, Z);
    input A1, A2, B;
    output Z;
endmodule
module OA21HVTD2 (A1, A2, B, Z);
    input A1, A2, B;
    output Z;
endmodule
module OA21HVTD4 (A1, A2, B, Z);
    input A1, A2, B;
    output Z;
endmodule
module OA221HVTD0 (A1, A2, B1, B2, C, Z);
    input A1, A2, B1, B2, C;
    output Z;
endmodule
module OA221HVTD1 (A1, A2, B1, B2, C, Z);
    input A1, A2, B1, B2, C;
    output Z;
endmodule
module OA221HVTD2 (A1, A2, B1, B2, C, Z);
    input A1, A2, B1, B2, C;
    output Z;
endmodule
module OA221HVTD4 (A1, A2, B1, B2, C, Z);
    input A1, A2, B1, B2, C;
    output Z;
endmodule
module OA222HVTD0 (A1, A2, B1, B2, C1, C2, Z);
    input A1, A2, B1, B2, C1, C2;
    output Z;
endmodule
module OA222HVTD1 (A1, A2, B1, B2, C1, C2, Z);
    input A1, A2, B1, B2, C1, C2;
    output Z;
endmodule
module OA222HVTD2 (A1, A2, B1, B2, C1, C2, Z);
    input A1, A2, B1, B2, C1, C2;
    output Z;
endmodule
module OA222HVTD4 (A1, A2, B1, B2, C1, C2, Z);
    input A1, A2, B1, B2, C1, C2;
    output Z;
endmodule
module OA22HVTD0 (A1, A2, B1, B2, Z);
    input A1, A2, B1, B2;
    output Z;
endmodule
module OA22HVTD1 (A1, A2, B1, B2, Z);
    input A1, A2, B1, B2;
    output Z;
endmodule
module OA22HVTD2 (A1, A2, B1, B2, Z);
    input A1, A2, B1, B2;
    output Z;
endmodule
module OA22HVTD4 (A1, A2, B1, B2, Z);
    input A1, A2, B1, B2;
    output Z;
endmodule
module OA31HVTD0 (A1, A2, A3, B, Z);
    input A1, A2, A3, B;
    output Z;
endmodule
module OA31HVTD1 (A1, A2, A3, B, Z);
    input A1, A2, A3, B;
    output Z;
endmodule
module OA31HVTD2 (A1, A2, A3, B, Z);
    input A1, A2, A3, B;
    output Z;
endmodule
module OA31HVTD4 (A1, A2, A3, B, Z);
    input A1, A2, A3, B;
    output Z;
endmodule
module OA32HVTD0 (A1, A2, A3, B1, B2, Z);
    input A1, A2, A3, B1, B2;
    output Z;
endmodule
module OA32HVTD1 (A1, A2, A3, B1, B2, Z);
    input A1, A2, A3, B1, B2;
    output Z;
endmodule
module OA32HVTD2 (A1, A2, A3, B1, B2, Z);
    input A1, A2, A3, B1, B2;
    output Z;
endmodule
module OA32HVTD4 (A1, A2, A3, B1, B2, Z);
    input A1, A2, A3, B1, B2;
    output Z;
endmodule
module OA33HVTD0 (A1, A2, A3, B1, B2, B3, Z);
    input A1, A2, A3, B1, B2, B3;
    output Z;
endmodule
module OA33HVTD1 (A1, A2, A3, B1, B2, B3, Z);
    input A1, A2, A3, B1, B2, B3;
    output Z;
endmodule
module OA33HVTD2 (A1, A2, A3, B1, B2, B3, Z);
    input A1, A2, A3, B1, B2, B3;
    output Z;
endmodule
module OA33HVTD4 (A1, A2, A3, B1, B2, B3, Z);
    input A1, A2, A3, B1, B2, B3;
    output Z;
endmodule
module OAI211HVTD0 (A1, A2, B, C, ZN);
    input A1, A2, B, C;
    output ZN;
endmodule
module OAI211HVTD1 (A1, A2, B, C, ZN);
    input A1, A2, B, C;
    output ZN;
endmodule
module OAI211HVTD2 (A1, A2, B, C, ZN);
    input A1, A2, B, C;
    output ZN;
endmodule
module OAI211HVTD4 (A1, A2, B, C, ZN);
    input A1, A2, B, C;
    output ZN;
endmodule
module OAI21HVTD0 (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
endmodule
module OAI21HVTD1 (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
endmodule
module OAI21HVTD2 (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
endmodule
module OAI21HVTD4 (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
endmodule
module OAI221HVTD0 (A1, A2, B1, B2, C, ZN);
    input A1, A2, B1, B2, C;
    output ZN;
endmodule
module OAI221HVTD1 (A1, A2, B1, B2, C, ZN);
    input A1, A2, B1, B2, C;
    output ZN;
endmodule
module OAI221HVTD2 (A1, A2, B1, B2, C, ZN);
    input A1, A2, B1, B2, C;
    output ZN;
endmodule
module OAI221HVTD4 (A1, A2, B1, B2, C, ZN);
    input A1, A2, B1, B2, C;
    output ZN;
endmodule
module OAI221XHVTD4 (A1, A2, B1, B2, C, ZN);
    input A1, A2, B1, B2, C;
    output ZN;
endmodule
module OAI222HVTD0 (A1, A2, B1, B2, C1, C2, ZN);
    input A1, A2, B1, B2, C1, C2;
    output ZN;
endmodule
module OAI222HVTD1 (A1, A2, B1, B2, C1, C2, ZN);
    input A1, A2, B1, B2, C1, C2;
    output ZN;
endmodule
module OAI222HVTD2 (A1, A2, B1, B2, C1, C2, ZN);
    input A1, A2, B1, B2, C1, C2;
    output ZN;
endmodule
module OAI222HVTD4 (A1, A2, B1, B2, C1, C2, ZN);
    input A1, A2, B1, B2, C1, C2;
    output ZN;
endmodule
module OAI222XHVTD4 (A1, A2, B1, B2, C1, C2, ZN);
    input A1, A2, B1, B2, C1, C2;
    output ZN;
endmodule
module OAI22HVTD0 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
endmodule
module OAI22HVTD1 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
endmodule
module OAI22HVTD2 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
endmodule
module OAI22HVTD4 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
endmodule
module OAI31HVTD0 (A1, A2, A3, B, ZN);
    input A1, A2, A3, B;
    output ZN;
endmodule
module OAI31HVTD1 (A1, A2, A3, B, ZN);
    input A1, A2, A3, B;
    output ZN;
endmodule
module OAI31HVTD2 (A1, A2, A3, B, ZN);
    input A1, A2, A3, B;
    output ZN;
endmodule
module OAI31HVTD4 (A1, A2, A3, B, ZN);
    input A1, A2, A3, B;
    output ZN;
endmodule
module OAI32HVTD0 (A1, A2, A3, B1, B2, ZN);
    input A1, A2, A3, B1, B2;
    output ZN;
endmodule
module OAI32HVTD1 (A1, A2, A3, B1, B2, ZN);
    input A1, A2, A3, B1, B2;
    output ZN;
endmodule
module OAI32HVTD2 (A1, A2, A3, B1, B2, ZN);
    input A1, A2, A3, B1, B2;
    output ZN;
endmodule
module OAI32HVTD4 (A1, A2, A3, B1, B2, ZN);
    input A1, A2, A3, B1, B2;
    output ZN;
endmodule
module OAI32XHVTD4 (A1, A2, A3, B1, B2, ZN);
    input A1, A2, A3, B1, B2;
    output ZN;
endmodule
module OAI33HVTD0 (A1, A2, A3, B1, B2, B3, ZN);
    input A1, A2, A3, B1, B2, B3;
    output ZN;
endmodule
module OAI33HVTD1 (A1, A2, A3, B1, B2, B3, ZN);
    input A1, A2, A3, B1, B2, B3;
    output ZN;
endmodule
module OAI33HVTD2 (A1, A2, A3, B1, B2, B3, ZN);
    input A1, A2, A3, B1, B2, B3;
    output ZN;
endmodule
module OAI33HVTD4 (A1, A2, A3, B1, B2, B3, ZN);
    input A1, A2, A3, B1, B2, B3;
    output ZN;
endmodule
module OAI33XHVTD4 (A1, A2, A3, B1, B2, B3, ZN);
    input A1, A2, A3, B1, B2, B3;
    output ZN;
endmodule
module OR2HVTD0 (A1, A2, Z);
    input A1, A2;
    output Z;
endmodule
module OR2HVTD1 (A1, A2, Z);
    input A1, A2;
    output Z;
endmodule
module OR2HVTD2 (A1, A2, Z);
    input A1, A2;
    output Z;
endmodule
module OR2HVTD4 (A1, A2, Z);
    input A1, A2;
    output Z;
endmodule
module OR2HVTD8 (A1, A2, Z);
    input A1, A2;
    output Z;
endmodule
module OR2XHVTD1 (A1, A2, Z);
    input A1, A2;
    output Z;
endmodule
module OR3HVTD0 (A1, A2, A3, Z);
    input A1, A2, A3;
    output Z;
endmodule
module OR3HVTD1 (A1, A2, A3, Z);
    input A1, A2, A3;
    output Z;
endmodule
module OR3HVTD2 (A1, A2, A3, Z);
    input A1, A2, A3;
    output Z;
endmodule
module OR3HVTD4 (A1, A2, A3, Z);
    input A1, A2, A3;
    output Z;
endmodule
module OR3HVTD8 (A1, A2, A3, Z);
    input A1, A2, A3;
    output Z;
endmodule
module OR3XHVTD1 (A1, A2, A3, Z);
    input A1, A2, A3;
    output Z;
endmodule
module OR4HVTD0 (A1, A2, A3, A4, Z);
    input A1, A2, A3, A4;
    output Z;
endmodule
module OR4HVTD1 (A1, A2, A3, A4, Z);
    input A1, A2, A3, A4;
    output Z;
endmodule
module OR4HVTD2 (A1, A2, A3, A4, Z);
    input A1, A2, A3, A4;
    output Z;
endmodule
module OR4HVTD4 (A1, A2, A3, A4, Z);
    input A1, A2, A3, A4;
    output Z;
endmodule
module OR4HVTD8 (A1, A2, A3, A4, Z);
    input A1, A2, A3, A4;
    output Z;
endmodule
module OR4XHVTD1 (A1, A2, A3, A4, Z);
    input A1, A2, A3, A4;
    output Z;
endmodule
module SDF4CQHVTD0 (SI, D, SE, CP, Q);
    input SI, D, SE, CP;
    output Q;
endmodule
module SDF4CQHVTD1 (SI, D, SE, CP, Q);
    input SI, D, SE, CP;
    output Q;
endmodule
module SDF4CQHVTD2 (SI, D, SE, CP, Q);
    input SI, D, SE, CP;
    output Q;
endmodule
module SDF4CQHVTD4 (SI, D, SE, CP, Q);
    input SI, D, SE, CP;
    output Q;
endmodule
module SDFCNHVTD0 (SI, D, SE, CP, CDN, Q, QN);
    input SI, D, SE, CP, CDN;
    output Q, QN;
endmodule
module SDFCNHVTD1 (SI, D, SE, CP, CDN, Q, QN);
    input SI, D, SE, CP, CDN;
    output Q, QN;
endmodule
module SDFCNHVTD2 (SI, D, SE, CP, CDN, Q, QN);
    input SI, D, SE, CP, CDN;
    output Q, QN;
endmodule
module SDFCNHVTD4 (SI, D, SE, CP, CDN, Q, QN);
    input SI, D, SE, CP, CDN;
    output Q, QN;
endmodule
module SDFCNQHVTD0 (SI, D, SE, CP, CDN, Q);
    input SI, D, SE, CP, CDN;
    output Q;
endmodule
module SDFCNQHVTD1 (SI, D, SE, CP, CDN, Q);
    input SI, D, SE, CP, CDN;
    output Q;
endmodule
module SDFCNQHVTD2 (SI, D, SE, CP, CDN, Q);
    input SI, D, SE, CP, CDN;
    output Q;
endmodule
module SDFCNQHVTD4 (SI, D, SE, CP, CDN, Q);
    input SI, D, SE, CP, CDN;
    output Q;
endmodule
module SDFCSNHVTD0 (SI, D, SE, CP, CDN, SDN, Q, QN);
    input SI, D, SE, CP, CDN, SDN;
    output Q, QN;
endmodule
module SDFCSNHVTD1 (SI, D, SE, CP, CDN, SDN, Q, QN);
    input SI, D, SE, CP, CDN, SDN;
    output Q, QN;
endmodule
module SDFCSNHVTD2 (SI, D, SE, CP, CDN, SDN, Q, QN);
    input SI, D, SE, CP, CDN, SDN;
    output Q, QN;
endmodule
module SDFCSNHVTD4 (SI, D, SE, CP, CDN, SDN, Q, QN);
    input SI, D, SE, CP, CDN, SDN;
    output Q, QN;
endmodule
module SDFCSNQHVTD0 (SI, D, SE, CP, CDN, SDN, Q);
    input SI, D, SE, CP, CDN, SDN;
    output Q;
endmodule
module SDFCSNQHVTD1 (SI, D, SE, CP, CDN, SDN, Q);
    input SI, D, SE, CP, CDN, SDN;
    output Q;
endmodule
module SDFCSNQHVTD2 (SI, D, SE, CP, CDN, SDN, Q);
    input SI, D, SE, CP, CDN, SDN;
    output Q;
endmodule
module SDFCSNQHVTD4 (SI, D, SE, CP, CDN, SDN, Q);
    input SI, D, SE, CP, CDN, SDN;
    output Q;
endmodule
module SDFHVTD0 (SI, D, SE, CP, Q, QN);
    input SI, D, SE, CP;
    output Q, QN;
endmodule
module SDFHVTD1 (SI, D, SE, CP, Q, QN);
    input SI, D, SE, CP;
    output Q, QN;
endmodule
module SDFHVTD2 (SI, D, SE, CP, Q, QN);
    input SI, D, SE, CP;
    output Q, QN;
endmodule
module SDFHVTD4 (SI, D, SE, CP, Q, QN);
    input SI, D, SE, CP;
    output Q, QN;
endmodule
module SDFKCNHVTD0 (SI, D, SE, CP, CN, Q, QN);
    input SI, D, SE, CP, CN;
    output Q, QN;
endmodule
module SDFKCNHVTD1 (SI, D, SE, CP, CN, Q, QN);
    input SI, D, SE, CP, CN;
    output Q, QN;
endmodule
module SDFKCNHVTD2 (SI, D, SE, CP, CN, Q, QN);
    input SI, D, SE, CP, CN;
    output Q, QN;
endmodule
module SDFKCNHVTD4 (SI, D, SE, CP, CN, Q, QN);
    input SI, D, SE, CP, CN;
    output Q, QN;
endmodule
module SDFKCNQHVTD0 (SI, D, SE, CP, CN, Q);
    input SI, D, SE, CP, CN;
    output Q;
endmodule
module SDFKCNQHVTD1 (SI, D, SE, CP, CN, Q);
    input SI, D, SE, CP, CN;
    output Q;
endmodule
module SDFKCNQHVTD2 (SI, D, SE, CP, CN, Q);
    input SI, D, SE, CP, CN;
    output Q;
endmodule
module SDFKCNQHVTD4 (SI, D, SE, CP, CN, Q);
    input SI, D, SE, CP, CN;
    output Q;
endmodule
module SDFKCSNHVTD0 (SI, D, SE, CP, CN, SN, Q, QN);
    input SI, D, SE, CP, CN, SN;
    output Q, QN;
endmodule
module SDFKCSNHVTD1 (SI, D, SE, CP, CN, SN, Q, QN);
    input SI, D, SE, CP, CN, SN;
    output Q, QN;
endmodule
module SDFKCSNHVTD2 (SI, D, SE, CP, CN, SN, Q, QN);
    input SI, D, SE, CP, CN, SN;
    output Q, QN;
endmodule
module SDFKCSNHVTD4 (SI, D, SE, CP, CN, SN, Q, QN);
    input SI, D, SE, CP, CN, SN;
    output Q, QN;
endmodule
module SDFKCSNQHVTD0 (SI, D, SE, CP, CN, SN, Q);
    input SI, D, SE, CP, CN, SN;
    output Q;
endmodule
module SDFKCSNQHVTD1 (SI, D, SE, CP, CN, SN, Q);
    input SI, D, SE, CP, CN, SN;
    output Q;
endmodule
module SDFKCSNQHVTD2 (SI, D, SE, CP, CN, SN, Q);
    input SI, D, SE, CP, CN, SN;
    output Q;
endmodule
module SDFKCSNQHVTD4 (SI, D, SE, CP, CN, SN, Q);
    input SI, D, SE, CP, CN, SN;
    output Q;
endmodule
module SDFKSNHVTD0 (SI, D, SE, CP, SN, Q, QN);
    input SI, D, SE, CP, SN;
    output Q, QN;
endmodule
module SDFKSNHVTD1 (SI, D, SE, CP, SN, Q, QN);
    input SI, D, SE, CP, SN;
    output Q, QN;
endmodule
module SDFKSNHVTD2 (SI, D, SE, CP, SN, Q, QN);
    input SI, D, SE, CP, SN;
    output Q, QN;
endmodule
module SDFKSNHVTD4 (SI, D, SE, CP, SN, Q, QN);
    input SI, D, SE, CP, SN;
    output Q, QN;
endmodule
module SDFKSNQHVTD0 (SI, D, SE, CP, SN, Q);
    input SI, D, SE, CP, SN;
    output Q;
endmodule
module SDFKSNQHVTD1 (SI, D, SE, CP, SN, Q);
    input SI, D, SE, CP, SN;
    output Q;
endmodule
module SDFKSNQHVTD2 (SI, D, SE, CP, SN, Q);
    input SI, D, SE, CP, SN;
    output Q;
endmodule
module SDFKSNQHVTD4 (SI, D, SE, CP, SN, Q);
    input SI, D, SE, CP, SN;
    output Q;
endmodule
module SDFNCNHVTD0 (SI, D, SE, CPN, CDN, Q, QN);
    input SI, D, SE, CPN, CDN;
    output Q, QN;
endmodule
module SDFNCNHVTD1 (SI, D, SE, CPN, CDN, Q, QN);
    input SI, D, SE, CPN, CDN;
    output Q, QN;
endmodule
module SDFNCNHVTD2 (SI, D, SE, CPN, CDN, Q, QN);
    input SI, D, SE, CPN, CDN;
    output Q, QN;
endmodule
module SDFNCNHVTD4 (SI, D, SE, CPN, CDN, Q, QN);
    input SI, D, SE, CPN, CDN;
    output Q, QN;
endmodule
module SDFNCSNHVTD0 (SI, D, SE, CPN, CDN, SDN, Q, QN);
    input SI, D, SE, CPN, CDN, SDN;
    output Q, QN;
endmodule
module SDFNCSNHVTD1 (SI, D, SE, CPN, CDN, SDN, Q, QN);
    input SI, D, SE, CPN, CDN, SDN;
    output Q, QN;
endmodule
module SDFNCSNHVTD2 (SI, D, SE, CPN, CDN, SDN, Q, QN);
    input SI, D, SE, CPN, CDN, SDN;
    output Q, QN;
endmodule
module SDFNCSNHVTD4 (SI, D, SE, CPN, CDN, SDN, Q, QN);
    input SI, D, SE, CPN, CDN, SDN;
    output Q, QN;
endmodule
module SDFNHVTD0 (SI, D, SE, CPN, Q, QN);
    input SI, D, SE, CPN;
    output Q, QN;
endmodule
module SDFNHVTD1 (SI, D, SE, CPN, Q, QN);
    input SI, D, SE, CPN;
    output Q, QN;
endmodule
module SDFNHVTD2 (SI, D, SE, CPN, Q, QN);
    input SI, D, SE, CPN;
    output Q, QN;
endmodule
module SDFNHVTD4 (SI, D, SE, CPN, Q, QN);
    input SI, D, SE, CPN;
    output Q, QN;
endmodule
module SDFNSNHVTD0 (SI, D, SE, CPN, SDN, Q, QN);
    input SI, D, SE, CPN, SDN;
    output Q, QN;
endmodule
module SDFNSNHVTD1 (SI, D, SE, CPN, SDN, Q, QN);
    input SI, D, SE, CPN, SDN;
    output Q, QN;
endmodule
module SDFNSNHVTD2 (SI, D, SE, CPN, SDN, Q, QN);
    input SI, D, SE, CPN, SDN;
    output Q, QN;
endmodule
module SDFNSNHVTD4 (SI, D, SE, CPN, SDN, Q, QN);
    input SI, D, SE, CPN, SDN;
    output Q, QN;
endmodule
module SDFQHVTD0 (SI, D, SE, CP, Q);
    input SI, D, SE, CP;
    output Q;
endmodule
module SDFQHVTD1 (SI, D, SE, CP, Q);
    input SI, D, SE, CP;
    output Q;
endmodule
module SDFQHVTD2 (SI, D, SE, CP, Q);
    input SI, D, SE, CP;
    output Q;
endmodule
module SDFQHVTD4 (SI, D, SE, CP, Q);
    input SI, D, SE, CP;
    output Q;
endmodule
module SDFQNHVTD0 (SI, D, SE, CP, QN);
    input SI, D, SE, CP;
    output QN;
endmodule
module SDFQNHVTD1 (SI, D, SE, CP, QN);
    input SI, D, SE, CP;
    output QN;
endmodule
module SDFQNHVTD2 (SI, D, SE, CP, QN);
    input SI, D, SE, CP;
    output QN;
endmodule
module SDFQNHVTD4 (SI, D, SE, CP, QN);
    input SI, D, SE, CP;
    output QN;
endmodule
module SDFSNHVTD0 (SI, D, SE, CP, SDN, Q, QN);
    input SI, D, SE, CP, SDN;
    output Q, QN;
endmodule
module SDFSNHVTD1 (SI, D, SE, CP, SDN, Q, QN);
    input SI, D, SE, CP, SDN;
    output Q, QN;
endmodule
module SDFSNHVTD2 (SI, D, SE, CP, SDN, Q, QN);
    input SI, D, SE, CP, SDN;
    output Q, QN;
endmodule
module SDFSNHVTD4 (SI, D, SE, CP, SDN, Q, QN);
    input SI, D, SE, CP, SDN;
    output Q, QN;
endmodule
module SDFSNQHVTD0 (SI, D, SE, CP, SDN, Q);
    input SI, D, SE, CP, SDN;
    output Q;
endmodule
module SDFSNQHVTD1 (SI, D, SE, CP, SDN, Q);
    input SI, D, SE, CP, SDN;
    output Q;
endmodule
module SDFSNQHVTD2 (SI, D, SE, CP, SDN, Q);
    input SI, D, SE, CP, SDN;
    output Q;
endmodule
module SDFSNQHVTD4 (SI, D, SE, CP, SDN, Q);
    input SI, D, SE, CP, SDN;
    output Q;
endmodule
module SDFXHVTD0 (DA, DB, SA, SI, SE, CP, Q, QN);
    input DA, DB, SA, SI, SE, CP;
    output Q, QN;
endmodule
module SDFXHVTD1 (DA, DB, SA, SI, SE, CP, Q, QN);
    input DA, DB, SA, SI, SE, CP;
    output Q, QN;
endmodule
module SDFXHVTD2 (DA, DB, SA, SI, SE, CP, Q, QN);
    input DA, DB, SA, SI, SE, CP;
    output Q, QN;
endmodule
module SDFXHVTD4 (DA, DB, SA, SI, SE, CP, Q, QN);
    input DA, DB, SA, SI, SE, CP;
    output Q, QN;
endmodule
module SDFXQHVTD0 (DA, DB, SA, SI, SE, CP, Q);
    input DA, DB, SA, SI, SE, CP;
    output Q;
endmodule
module SDFXQHVTD1 (DA, DB, SA, SI, SE, CP, Q);
    input DA, DB, SA, SI, SE, CP;
    output Q;
endmodule
module SDFXQHVTD2 (DA, DB, SA, SI, SE, CP, Q);
    input DA, DB, SA, SI, SE, CP;
    output Q;
endmodule
module SDFXQHVTD4 (DA, DB, SA, SI, SE, CP, Q);
    input DA, DB, SA, SI, SE, CP;
    output Q;
endmodule
module SEDF4CQHVTD0 (E, SE, CP, SI, D, Q);
    input E, SE, CP, SI, D; 
    output Q;
endmodule
module SEDF4CQHVTD1 (E, SE, CP, SI, D, Q);
    input E, SE, CP, SI, D; 
    output Q;
endmodule
module SEDF4CQHVTD2 (E, SE, CP, SI, D, Q);
    input E, SE, CP, SI, D; 
    output Q;
endmodule
module SEDF4CQHVTD4 (E, SE, CP, SI, D, Q);
    input E, SE, CP, SI, D; 
    output Q;
endmodule
module SEDFCNHVTD0 (E, SE, CP, SI, D, CDN, Q, QN);
    input E, SE, CP, SI, D, CDN; 
    output Q, QN;
endmodule
module SEDFCNHVTD1 (E, SE, CP, SI, D, CDN, Q, QN);
    input E, SE, CP, SI, D, CDN; 
    output Q, QN;
endmodule
module SEDFCNHVTD2 (E, SE, CP, SI, D, CDN, Q, QN);
    input E, SE, CP, SI, D, CDN; 
    output Q, QN;
endmodule
module SEDFCNHVTD4 (E, SE, CP, SI, D, CDN, Q, QN);
    input E, SE, CP, SI, D, CDN; 
    output Q, QN;
endmodule
module SEDFCNQHVTD0 (E, SE, CP, SI, D, CDN, Q);
    input E, SE, CP, SI, D, CDN; 
    output Q;
endmodule
module SEDFCNQHVTD1 (E, SE, CP, SI, D, CDN, Q);
    input E, SE, CP, SI, D, CDN; 
    output Q;
endmodule
module SEDFCNQHVTD2 (E, SE, CP, SI, D, CDN, Q);
    input E, SE, CP, SI, D, CDN; 
    output Q;
endmodule
module SEDFCNQHVTD4 (E, SE, CP, SI, D, CDN, Q);
    input E, SE, CP, SI, D, CDN; 
    output Q;
endmodule
module SEDFHVTD0 (E, SE, CP, SI, D, Q, QN);
    input E, SE, CP, SI, D; 
    output Q, QN;
endmodule
module SEDFHVTD1 (E, SE, CP, SI, D, Q, QN);
    input E, SE, CP, SI, D; 
    output Q, QN;
endmodule
module SEDFHVTD2 (E, SE, CP, SI, D, Q, QN);
    input E, SE, CP, SI, D; 
    output Q, QN;
endmodule
module SEDFHVTD4 (E, SE, CP, SI, D, Q, QN);
    input E, SE, CP, SI, D; 
    output Q, QN;
endmodule
module SEDFKCNHVTD0 (SI, D, E, SE, CP, CN, Q, QN);
    input SI, D, SE, CP, CN, E;
    output Q, QN;
endmodule
module SEDFKCNHVTD1 (SI, D, E, SE, CP, CN, Q, QN);
    input SI, D, SE, CP, CN, E;
    output Q, QN;
endmodule
module SEDFKCNHVTD2 (SI, D, E, SE, CP, CN, Q, QN);
    input SI, D, SE, CP, CN, E;
    output Q, QN;
endmodule
module SEDFKCNHVTD4 (SI, D, E, SE, CP, CN, Q, QN);
    input SI, D, SE, CP, CN, E;
    output Q, QN;
endmodule
module SEDFKCNQHVTD0 (SI, D, E, SE, CP, CN, Q);
    input SI, D, SE, CP, CN, E;
    output Q;
endmodule
module SEDFKCNQHVTD1 (SI, D, E, SE, CP, CN, Q);
    input SI, D, SE, CP, CN, E;
    output Q;
endmodule
module SEDFKCNQHVTD2 (SI, D, E, SE, CP, CN, Q);
    input SI, D, SE, CP, CN, E;
    output Q;
endmodule
module SEDFKCNQHVTD4 (SI, D, E, SE, CP, CN, Q);
    input SI, D, SE, CP, CN, E;
    output Q;
endmodule
module SEDFQHVTD0 (E, SE, CP, SI, D, Q);
    input E, SE, CP, SI, D; 
    output Q;
endmodule
module SEDFQHVTD1 (E, SE, CP, SI, D, Q);
    input E, SE, CP, SI, D; 
    output Q;
endmodule
module SEDFQHVTD2 (E, SE, CP, SI, D, Q);
    input E, SE, CP, SI, D; 
    output Q;
endmodule
module SEDFQHVTD4 (E, SE, CP, SI, D, Q);
    input E, SE, CP, SI, D; 
    output Q;
endmodule
module SEDFQNHVTD0 (E, SE, CP, SI, D, QN);
    input E, SE, CP, SI, D; 
    output QN;
endmodule
module SEDFQNHVTD1 (E, SE, CP, SI, D, QN);
    input E, SE, CP, SI, D; 
    output QN;
endmodule
module SEDFQNHVTD2 (E, SE, CP, SI, D, QN);
    input E, SE, CP, SI, D; 
    output QN;
endmodule
module SEDFQNHVTD4 (E, SE, CP, SI, D, QN);
    input E, SE, CP, SI, D; 
    output QN;
endmodule
module TIEHHVT (Z);
  output  Z;
endmodule
module TIELHVT (ZN);
  output  ZN;
endmodule
module XNR2HVTD0 (A1, A2, ZN);
  input		A1, A2;
  output 	ZN;
endmodule
module XNR2HVTD1 (A1, A2, ZN);
  input		A1, A2;
  output 	ZN;
endmodule
module XNR2HVTD2 (A1, A2, ZN);
  input		A1, A2;
  output 	ZN;
endmodule
module XNR2HVTD4 (A1, A2, ZN);
  input		A1, A2;
  output 	ZN;
endmodule
module XNR3HVTD0 (A1, A2, A3, ZN);
  input A1, A2, A3;
  output ZN;
endmodule
module XNR3HVTD1 (A1, A2, A3, ZN);
  input A1, A2, A3;
  output ZN;
endmodule
module XNR3HVTD2 (A1, A2, A3, ZN);
  input A1, A2, A3;
  output ZN;
endmodule
module XNR3HVTD4 (A1, A2, A3, ZN);
  input A1, A2, A3;
  output ZN;
endmodule
module XNR4HVTD0 (A1, A2, A3, A4, ZN);
  input 	A1, A2, A3, A4;
  output 	ZN;
endmodule
module XNR4HVTD1 (A1, A2, A3, A4, ZN);
  input 	A1, A2, A3, A4;
  output 	ZN;
endmodule
module XNR4HVTD2 (A1, A2, A3, A4, ZN);
  input 	A1, A2, A3, A4;
  output 	ZN;
endmodule
module XNR4HVTD4 (A1, A2, A3, A4, ZN);
  input 	A1, A2, A3, A4;
  output 	ZN;
endmodule
module XOR2HVTD0 (A1, A2, Z);
  input 	A1, A2;
  output 	Z;
endmodule
module XOR2HVTD1 (A1, A2, Z);
  input 	A1, A2;
  output 	Z;
endmodule
module XOR2HVTD2 (A1, A2, Z);
  input 	A1, A2;
  output 	Z;
endmodule
module XOR2HVTD4 (A1, A2, Z);
  input 	A1, A2;
  output 	Z;
endmodule
module XOR3HVTD0 (A1, A2, A3, Z);
  input A1, A2, A3;
  output Z;
endmodule
module XOR3HVTD1 (A1, A2, A3, Z);
  input A1, A2, A3;
  output Z;
endmodule
module XOR3HVTD2 (A1, A2, A3, Z);
  input A1, A2, A3;
  output Z;
endmodule
module XOR3HVTD4 (A1, A2, A3, Z);
  input A1, A2, A3;
  output Z;
endmodule
module XOR4HVTD0 (A1, A2, A3, A4, Z);
  input 	A1, A2, A3, A4;
  output 	Z;
endmodule
module XOR4HVTD1 (A1, A2, A3, A4, Z);
  input 	A1, A2, A3, A4;
  output 	Z;
endmodule
module XOR4HVTD2 (A1, A2, A3, A4, Z);
  input 	A1, A2, A3, A4;
  output 	Z;
endmodule
module XOR4HVTD4 (A1, A2, A3, A4, Z);
  input 	A1, A2, A3, A4;
  output 	Z;
endmodule
