module invalidSyntax;
  reg test
endmodule
