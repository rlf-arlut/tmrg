module invalidSyntax;
  reg2 test;
endmodule
