
module top (output E1A);
  // tmrg default triplicate
  mod d0 (.E1(E1A));
endmodule

module mod (output E1);
// tmrg default triplicate
endmodule

