module wireTest;
  // tmrg do_not_triplicate i
  // tmrg triplicate j
  wire i,j;
endmodule
