module comb01( 
  input [7:0]  in1, 
  out2,
  output [P:2] dd,
  inout [X:D] pp
  );
  output [1:2] out5, x2;
  output x,y;
  input [1:2] out5,x2;

  assign out= #1 fun(in)
  +in2,out2=i1+in2;
  assign out4=fun(in)+in2, out3=i1+in2;
  always @(in1)
  begin
    out1=in1;
    out1=in1;
    i2<=in1;
    if (in) 
      x<=2'b0;
    if (x && y==1'b1) 
      a=0;
    else
      begin
        v=2;
        if (d) begin y=2; end
      end
  end

  always
    out1=in1;
  
  modulename inst1 (.d(s)) , inst2 (.d(s) , ds );
endmodule

