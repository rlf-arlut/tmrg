module vote01 (in,out);
  // tmrg default triplicate
  input in;
  output out;
  wire inVoted = in;
  assign out = inVoted;
endmodule
