module b;
    reg [1:0] x = 5'd3;
endmodule
