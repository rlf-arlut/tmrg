module divider(
  input clkin,
  output clkout1,
  output clkout2
);

  // tmrg default triplicate
  // tmrg do_not_triplicate clkout2

endmodule
