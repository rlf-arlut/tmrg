module real_test(
  input real i,
  output real o
);
  assign o = i;
endmodule
