`resetall
module wiretest(input clk,input d, output q);
wire [7:0] re[0:1],r5;
wire [7:0] registers2,r3,r4;
reg [7:0] registers3[0:13];

endmodule
