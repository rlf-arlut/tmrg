module m1();
endmodule
module m2();
endmodule
