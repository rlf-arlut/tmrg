module test;
localparam W=9;
localparam H=2;
integer i=0;
integer k=9,j=1;
integer kk=W-H;
integer maxWH=(W>H)?W:H;
integer absWH=(W>H)?W-H:H-W;
endmodule
