module m3(i,o);
input i;
output o;
/* xxx instXXX(.i(i),.o(o)); */
endmodule

