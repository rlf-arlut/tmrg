module comb01( 
  input [7:0]  in, 
  input [7:0]  in2, 
  output [8:0] out
  );
  assign out=in+in2;

endmodule
