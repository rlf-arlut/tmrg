`include "always.v"
module x;
wire clk,d,q;
al alinst(.clk(clk),.d(d),.q(q));
endmodule

// _tmrg include.v -vv  --include --inc-dir="."
