module test;
  function static integer mux;
    input a, b, c, d;
  endfunction
endmodule

