module package_import;
  import my_package_pkg::ZERO;
  import my_package_pkg::ONE, my_package_pkg::TWO;
  import my_package_pkg::*;
endmodule
