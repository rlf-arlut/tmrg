module AN2D0 (A1, A2, Z);
    input A1, A2;
    output Z;
endmodule
module AN2D1 (A1, A2, Z);
    input A1, A2;
    output Z;
endmodule
module AN2D2 (A1, A2, Z);
    input A1, A2;
    output Z;
endmodule
module AN2D4 (A1, A2, Z);
    input A1, A2;
    output Z;
endmodule
module AN2D8 (A1, A2, Z);
    input A1, A2;
    output Z;
endmodule
module AN2XD1 (A1, A2, Z);
    input A1, A2;
    output Z;
endmodule
module AN3D0 (A1, A2, A3, Z);
    input A1, A2, A3;
    output Z;
endmodule
module AN3D1 (A1, A2, A3, Z);
    input A1, A2, A3;
    output Z;
endmodule
module AN3D2 (A1, A2, A3, Z);
    input A1, A2, A3;
    output Z;
endmodule
module AN3D4 (A1, A2, A3, Z);
    input A1, A2, A3;
    output Z;
endmodule
module AN3D8 (A1, A2, A3, Z);
    input A1, A2, A3;
    output Z;
endmodule
module AN3XD1 (A1, A2, A3, Z);
    input A1, A2, A3;
    output Z;
endmodule
module AN4D0 (A1, A2, A3, A4, Z);
    input A1, A2, A3, A4;
    output Z;
endmodule
module AN4D1 (A1, A2, A3, A4, Z);
    input A1, A2, A3, A4;
    output Z;
endmodule
module AN4D2 (A1, A2, A3, A4, Z);
    input A1, A2, A3, A4;
    output Z;
endmodule
module AN4D4 (A1, A2, A3, A4, Z);
    input A1, A2, A3, A4;
    output Z;
endmodule
module AN4D8 (A1, A2, A3, A4, Z);
    input A1, A2, A3, A4;
    output Z;
endmodule
module AN4XD1 (A1, A2, A3, A4, Z);
    input A1, A2, A3, A4;
    output Z;
endmodule
module ANTENNA (I);
  input I;
endmodule
module AO211D0 (A1, A2, B, C, Z);
    input A1, A2, B, C;
    output Z;
endmodule
module AO211D1 (A1, A2, B, C, Z);
    input A1, A2, B, C;
    output Z;
endmodule
module AO211D2 (A1, A2, B, C, Z);
    input A1, A2, B, C;
    output Z;
endmodule
module AO211D4 (A1, A2, B, C, Z);
    input A1, A2, B, C;
    output Z;
endmodule
module AO21D0 (A1, A2, B, Z);
    input A1, A2, B;
    output Z;
endmodule
module AO21D1 (A1, A2, B, Z);
    input A1, A2, B;
    output Z;
endmodule
module AO21D2 (A1, A2, B, Z);
    input A1, A2, B;
    output Z;
endmodule
module AO21D4 (A1, A2, B, Z);
    input A1, A2, B;
    output Z;
endmodule
module AO221D0 (A1, A2, B1, B2, C, Z);
    input A1, A2, B1, B2, C;
    output Z;
endmodule
module AO221D1 (A1, A2, B1, B2, C, Z);
    input A1, A2, B1, B2, C;
    output Z;
endmodule
module AO221D2 (A1, A2, B1, B2, C, Z);
    input A1, A2, B1, B2, C;
    output Z;
endmodule
module AO221D4 (A1, A2, B1, B2, C, Z);
    input A1, A2, B1, B2, C;
    output Z;
endmodule
module AO222D0 (A1, A2, B1, B2, C1, C2, Z);
    input A1, A2, B1, B2, C1, C2;
    output Z;
endmodule
module AO222D1 (A1, A2, B1, B2, C1, C2, Z);
    input A1, A2, B1, B2, C1, C2;
    output Z;
endmodule
module AO222D2 (A1, A2, B1, B2, C1, C2, Z);
    input A1, A2, B1, B2, C1, C2;
    output Z;
endmodule
module AO222D4 (A1, A2, B1, B2, C1, C2, Z);
    input A1, A2, B1, B2, C1, C2;
    output Z;
endmodule
module AO22D0 (A1, A2, B1, B2, Z);
    input A1, A2, B1, B2;
    output Z;
endmodule
module AO22D1 (A1, A2, B1, B2, Z);
    input A1, A2, B1, B2;
    output Z;
endmodule
module AO22D2 (A1, A2, B1, B2, Z);
    input A1, A2, B1, B2;
    output Z;
endmodule
module AO22D4 (A1, A2, B1, B2, Z);
    input A1, A2, B1, B2;
    output Z;
endmodule
module AO31D0 (A1, A2, A3, B, Z);
    input A1, A2, A3, B;
    output Z;
endmodule
module AO31D1 (A1, A2, A3, B, Z);
    input A1, A2, A3, B;
    output Z;
endmodule
module AO31D2 (A1, A2, A3, B, Z);
    input A1, A2, A3, B;
    output Z;
endmodule
module AO31D4 (A1, A2, A3, B, Z);
    input A1, A2, A3, B;
    output Z;
endmodule
module AO32D0 (A1, A2, A3, B1, B2, Z);
    input A1, A2, A3, B1, B2;
    output Z;
endmodule
module AO32D1 (A1, A2, A3, B1, B2, Z);
    input A1, A2, A3, B1, B2;
    output Z;
endmodule
module AO32D2 (A1, A2, A3, B1, B2, Z);
    input A1, A2, A3, B1, B2;
    output Z;
endmodule
module AO32D4 (A1, A2, A3, B1, B2, Z);
    input A1, A2, A3, B1, B2;
    output Z;
endmodule
module AO33D0 (A1, A2, A3, B1, B2, B3, Z);
    input A1, A2, A3, B1, B2, B3;
    output Z;
endmodule
module AO33D1 (A1, A2, A3, B1, B2, B3, Z);
    input A1, A2, A3, B1, B2, B3;
    output Z;
endmodule
module AO33D2 (A1, A2, A3, B1, B2, B3, Z);
    input A1, A2, A3, B1, B2, B3;
    output Z;
endmodule
module AO33D4 (A1, A2, A3, B1, B2, B3, Z);
    input A1, A2, A3, B1, B2, B3;
    output Z;
endmodule
module AOI211D0 (A1, A2, B, C, ZN);
    input A1, A2, B, C;
    output ZN;
endmodule
module AOI211D1 (A1, A2, B, C, ZN);
    input A1, A2, B, C;
    output ZN;
endmodule
module AOI211D2 (A1, A2, B, C, ZN);
    input A1, A2, B, C;
    output ZN;
endmodule
module AOI211D4 (A1, A2, B, C, ZN);
    input A1, A2, B, C;
    output ZN;
endmodule
module AOI211XD0 (A1, A2, B, C, ZN);
    input A1, A2, B, C;
    output ZN;
endmodule
module AOI211XD1 (A1, A2, B, C, ZN);
    input A1, A2, B, C;
    output ZN;
endmodule
module AOI211XD2 (A1, A2, B, C, ZN);
    input A1, A2, B, C;
    output ZN;
endmodule
module AOI211XD4 (A1, A2, B, C, ZN);
    input A1, A2, B, C;
    output ZN;
endmodule
module AOI21D0 (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
endmodule
module AOI21D1 (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
endmodule
module AOI21D2 (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
endmodule
module AOI21D4 (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
endmodule
module AOI221D0 (A1, A2, B1, B2, C, ZN);
    input A1, A2, B1, B2, C;
    output ZN;
endmodule
module AOI221D1 (A1, A2, B1, B2, C, ZN);
    input A1, A2, B1, B2, C;
    output ZN;
endmodule
module AOI221D2 (A1, A2, B1, B2, C, ZN);
    input A1, A2, B1, B2, C;
    output ZN;
endmodule
module AOI221D4 (A1, A2, B1, B2, C, ZN);
    input A1, A2, B1, B2, C;
    output ZN;
endmodule
module AOI221XD4 (A1, A2, B1, B2, C, ZN);
    input A1, A2, B1, B2, C;
    output ZN;
endmodule
module AOI222D0 (A1, A2, B1, B2, C1, C2, ZN);
    input A1, A2, B1, B2, C1, C2;
    output ZN;
endmodule
module AOI222D1 (A1, A2, B1, B2, C1, C2, ZN);
    input A1, A2, B1, B2, C1, C2;
    output ZN;
endmodule
module AOI222D2 (A1, A2, B1, B2, C1, C2, ZN);
    input A1, A2, B1, B2, C1, C2;
    output ZN;
endmodule
module AOI222D4 (A1, A2, B1, B2, C1, C2, ZN);
    input A1, A2, B1, B2, C1, C2;
    output ZN;
endmodule
module AOI222XD4 (A1, A2, B1, B2, C1, C2, ZN);
    input A1, A2, B1, B2, C1, C2;
    output ZN;
endmodule
module AOI22D0 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
endmodule
module AOI22D1 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
endmodule
module AOI22D2 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
endmodule
module AOI22D4 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
endmodule
module AOI31D0 (A1, A2, A3, B, ZN);
    input A1, A2, A3, B;
    output ZN;
endmodule
module AOI31D1 (A1, A2, A3, B, ZN);
    input A1, A2, A3, B;
    output ZN;
endmodule
module AOI31D2 (A1, A2, A3, B, ZN);
    input A1, A2, A3, B;
    output ZN;
endmodule
module AOI31D4 (A1, A2, A3, B, ZN);
    input A1, A2, A3, B;
    output ZN;
endmodule
module AOI32D0 (A1, A2, A3, B1, B2, ZN);
    input A1, A2, A3, B1, B2;
    output ZN;
endmodule
module AOI32D1 (A1, A2, A3, B1, B2, ZN);
    input A1, A2, A3, B1, B2;
    output ZN;
endmodule
module AOI32D2 (A1, A2, A3, B1, B2, ZN);
    input A1, A2, A3, B1, B2;
    output ZN;
endmodule
module AOI32D4 (A1, A2, A3, B1, B2, ZN);
    input A1, A2, A3, B1, B2;
    output ZN;
endmodule
module AOI32XD4 (A1, A2, A3, B1, B2, ZN);
    input A1, A2, A3, B1, B2;
    output ZN;
endmodule
module AOI33D0 (A1, A2, A3, B1, B2, B3, ZN);
    input A1, A2, A3, B1, B2, B3;
    output ZN;
endmodule
module AOI33D1 (A1, A2, A3, B1, B2, B3, ZN);
    input A1, A2, A3, B1, B2, B3;
    output ZN;
endmodule
module AOI33D2 (A1, A2, A3, B1, B2, B3, ZN);
    input A1, A2, A3, B1, B2, B3;
    output ZN;
endmodule
module AOI33D4 (A1, A2, A3, B1, B2, B3, ZN);
    input A1, A2, A3, B1, B2, B3;
    output ZN;
endmodule
module AOI33XD4 (A1, A2, A3, B1, B2, B3, ZN);
    input A1, A2, A3, B1, B2, B3;
    output ZN;
endmodule
module BENCD1 (M0, M1, M2, X2, A, S);
    input M0, M1, M2;
    output X2, A, S;
endmodule
module BENCD2 (M0, M1, M2, X2, A, S);
    input M0, M1, M2;
    output X2, A, S;
endmodule
module BENCD4 (M0, M1, M2, X2, A, S);
    input M0, M1, M2;
    output X2, A, S;
endmodule
module BMLD1 (X2, A, S, M0, M1, PP);
  input		X2, A, S, M0, M1;
  output	PP;
endmodule
module BMLD2 (X2, A, S, M0, M1, PP);
  input		X2, A, S, M0, M1;
  output	PP;
endmodule
module BMLD4 (X2, A, S, M0, M1, PP);
  input		X2, A, S, M0, M1;
  output	PP;
endmodule
module BUFFD0 (I, Z);
    input I;
    output Z;
endmodule
module BUFFD1 (I, Z);
    input I;
    output Z;
endmodule
module BUFFD12 (I, Z);
    input I;
    output Z;
endmodule
module BUFFD16 (I, Z);
    input I;
    output Z;
endmodule
module BUFFD2 (I, Z);
    input I;
    output Z;
endmodule
module BUFFD20 (I, Z);
    input I;
    output Z;
endmodule
module BUFFD24 (I, Z);
    input I;
    output Z;
endmodule
module BUFFD3 (I, Z);
    input I;
    output Z;
endmodule
module BUFFD4 (I, Z);
    input I;
    output Z;
endmodule
module BUFFD6 (I, Z);
    input I;
    output Z;
endmodule
module BUFFD8 (I, Z);
    input I;
    output Z;
endmodule
module BUFTD0 (I, OE, Z);
    input I, OE;
    output Z;
endmodule
module BUFTD1 (I, OE, Z);
    input I, OE;
    output Z;
endmodule
module BUFTD12 (I, OE, Z);
    input I, OE;
    output Z;
endmodule
module BUFTD16 (I, OE, Z);
    input I, OE;
    output Z;
endmodule
module BUFTD2 (I, OE, Z);
    input I, OE;
    output Z;
endmodule
module BUFTD20 (I, OE, Z);
    input I, OE;
    output Z;
endmodule
module BUFTD24 (I, OE, Z);
    input I, OE;
    output Z;
endmodule
module BUFTD3 (I, OE, Z);
    input I, OE;
    output Z;
endmodule
module BUFTD4 (I, OE, Z);
    input I, OE;
    output Z;
endmodule
module BUFTD6 (I, OE, Z);
    input I, OE;
    output Z;
endmodule
module BUFTD8 (I, OE, Z);
    input I, OE;
    output Z;
endmodule
module CKAN2D0 (A1, A2, Z);
    input A1, A2;
    output Z;
endmodule
module CKAN2D1 (A1, A2, Z);
    input A1, A2;
    output Z;
endmodule
module CKAN2D2 (A1, A2, Z);
    input A1, A2;
    output Z;
endmodule
module CKAN2D4 (A1, A2, Z);
    input A1, A2;
    output Z;
endmodule
module CKAN2D8 (A1, A2, Z);
    input A1, A2;
    output Z;
endmodule
module CKBD0 (I, Z);
    input I;
    output Z;
endmodule
module CKBD1 (I, Z);
    input I;
    output Z;
endmodule
module CKBD12 (I, Z);
    input I;
    output Z;
endmodule
module CKBD16 (I, Z);
    input I;
    output Z;
endmodule
module CKBD2 (I, Z);
    input I;
    output Z;
endmodule
module CKBD20 (I, Z);
    input I;
    output Z;
endmodule
module CKBD24 (I, Z);
    input I;
    output Z;
endmodule
module CKBD3 (I, Z);
    input I;
    output Z;
endmodule
module CKBD4 (I, Z);
    input I;
    output Z;
endmodule
module CKBD6 (I, Z);
    input I;
    output Z;
endmodule
module CKBD8 (I, Z);
    input I;
    output Z;
endmodule
module CKLHQD1 ( Q, TE, CPN, E );
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input TE, CPN, E;
    output Q;
endmodule
module CKLHQD12 ( Q, TE, CPN, E );
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input TE, CPN, E;
    output Q;
endmodule
module CKLHQD16 ( Q, TE, CPN, E );
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input TE, CPN, E;
    output Q;
endmodule
module CKLHQD2 ( Q, TE, CPN, E );
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input TE, CPN, E;
    output Q;
endmodule
module CKLHQD20 ( Q, TE, CPN, E );
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input TE, CPN, E;
    output Q;
endmodule
module CKLHQD24 ( Q, TE, CPN, E );
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input TE, CPN, E;
    output Q;
endmodule
module CKLHQD3 ( Q, TE, CPN, E );
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input TE, CPN, E;
    output Q;
endmodule
module CKLHQD4 ( Q, TE, CPN, E );
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input TE, CPN, E;
    output Q;
endmodule
module CKLHQD6 ( Q, TE, CPN, E );
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input TE, CPN, E;
    output Q;
endmodule
module CKLHQD8 ( Q, TE, CPN, E );
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input TE, CPN, E;
    output Q;
endmodule
module CKLNQD1 (TE, E, CP, Q);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input TE, E, CP;
    output Q;
endmodule
module CKLNQD12 (TE, E, CP, Q);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input TE, E, CP;
    output Q;
endmodule
module CKLNQD16 (TE, E, CP, Q);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input TE, E, CP;
    output Q;
endmodule
module CKLNQD2 (TE, E, CP, Q);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input TE, E, CP;
    output Q;
endmodule
module CKLNQD20 (TE, E, CP, Q);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input TE, E, CP;
    output Q;
endmodule
module CKLNQD24 (TE, E, CP, Q);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input TE, E, CP;
    output Q;
endmodule
module CKLNQD3 (TE, E, CP, Q);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input TE, E, CP;
    output Q;
endmodule
module CKLNQD4 (TE, E, CP, Q);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input TE, E, CP;
    output Q;
endmodule
module CKLNQD6 (TE, E, CP, Q);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input TE, E, CP;
    output Q;
endmodule
module CKLNQD8 (TE, E, CP, Q);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input TE, E, CP;
    output Q;
endmodule
module CKMUX2D0 (I0, I1, S, Z);
  input		I0, I1, S;
  output	Z;
endmodule
module CKMUX2D1 (I0, I1, S, Z);
  input		I0, I1, S;
  output	Z;
endmodule
module CKMUX2D2 (I0, I1, S, Z);
  input		I0, I1, S;
  output	Z;
endmodule
module CKMUX2D4 (I0, I1, S, Z);
  input		I0, I1, S;
  output	Z;
endmodule
module CKND0 (I, ZN);
    input I;
    output ZN;
endmodule
module CKND1 (I, ZN);
    input I;
    output ZN;
endmodule
module CKND12 (I, ZN);
    input I;
    output ZN;
endmodule
module CKND16 (I, ZN);
    input I;
    output ZN;
endmodule
module CKND2 (I, ZN);
    input I;
    output ZN;
endmodule
module CKND20 (I, ZN);
    input I;
    output ZN;
endmodule
module CKND24 (I, ZN);
    input I;
    output ZN;
endmodule
module CKND2D0 (A1, A2, ZN);
    input A1, A2;
    output ZN;
endmodule
module CKND2D1 (A1, A2, ZN);
    input A1, A2;
    output ZN;
endmodule
module CKND2D2 (A1, A2, ZN);
    input A1, A2;
    output ZN;
endmodule
module CKND2D3 (A1, A2, ZN);
    input A1, A2;
    output ZN;
endmodule
module CKND2D4 (A1, A2, ZN);
    input A1, A2;
    output ZN;
endmodule
module CKND2D8 (A1, A2, ZN);
    input A1, A2;
    output ZN;
endmodule
module CKND3 (I, ZN);
    input I;
    output ZN;
endmodule
module CKND4 (I, ZN);
    input I;
    output ZN;
endmodule
module CKND6 (I, ZN);
    input I;
    output ZN;
endmodule
module CKND8 (I, ZN);
    input I;
    output ZN;
endmodule
module CKXOR2D0 (A1, A2, Z);
  input 	A1, A2;
  output 	Z;
endmodule
module CKXOR2D1 (A1, A2, Z);
  input 	A1, A2;
  output 	Z;
endmodule
module CKXOR2D2 (A1, A2, Z);
  input 	A1, A2;
  output 	Z;
endmodule
module CKXOR2D4 (A1, A2, Z);
  input 	A1, A2;
  output 	Z;
endmodule
module CMPE42D1 (A, B, C, D, CIX, S, COX, CO);
input A, B, C, D, CIX;
output S, COX, CO;
endmodule
module CMPE42D2 (A, B, C, D, CIX, S, COX, CO);
input A, B, C, D, CIX;
output S, COX, CO;
endmodule
module DCAP;
endmodule
module DCAP16;
endmodule
module DCAP32;
endmodule
module DCAP4;
endmodule
module DCAP64;
endmodule
module DCAP8;
endmodule
module DEL0 (I, Z);
    input I;
    output Z;
endmodule
module DEL005 (I, Z);
    input I;
    output Z;
endmodule
module DEL01 (I, Z);
    input I;
    output Z;
endmodule
module DEL015 (I, Z);
    input I;
    output Z;
endmodule
module DEL02 (I, Z);
    input I;
    output Z;
endmodule
module DEL1 (I, Z);
    input I;
    output Z;
endmodule
module DEL2 (I, Z);
    input I;
    output Z;
endmodule
module DEL3 (I, Z);
    input I;
    output Z;
endmodule
module DEL4 (I, Z);
    input I;
    output Z;
endmodule
module DFCND1 (D, CP, CDN, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input D, CP, CDN;
    output Q, QN;
endmodule
module DFCND2 (D, CP, CDN, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input D, CP, CDN;
    output Q, QN;
endmodule
module DFCND4 (D, CP, CDN, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input D, CP, CDN;
    output Q, QN;
endmodule
module DFCNQD1 (D, CP, CDN, Q);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input D, CP, CDN;
    output Q;
endmodule
module DFCNQD2 (D, CP, CDN, Q);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input D, CP, CDN;
    output Q;
endmodule
module DFCNQD4 (D, CP, CDN, Q);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input D, CP, CDN;
    output Q;
endmodule
module DFCSND1 (D, CP, CDN, SDN, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input D, CP, CDN, SDN;
    output Q, QN;
endmodule
module DFCSND2 (D, CP, CDN, SDN, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input D, CP, CDN, SDN;
    output Q, QN;
endmodule
module DFCSND4 (D, CP, CDN, SDN, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input D, CP, CDN, SDN;
    output Q, QN;
endmodule
module DFCSNQD1 (D, CP, CDN, SDN, Q);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input D, CP, CDN, SDN;
    output Q;
endmodule
module DFCSNQD2 (D, CP, CDN, SDN, Q);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input D, CP, CDN, SDN;
    output Q;
endmodule
module DFCSNQD4 (D, CP, CDN, SDN, Q);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input D, CP, CDN, SDN;
    output Q;
endmodule
module DFD1 (D, CP, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input D, CP;
    output Q, QN;
endmodule
module DFD2 (D, CP, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input D, CP;
    output Q, QN;
endmodule
module DFD4 (D, CP, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input D, CP;
    output Q, QN;
endmodule
module DFKCND1 (D, CP, CN, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input D, CP, CN;
    output Q, QN;
endmodule
module DFKCND2 (D, CP, CN, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input D, CP, CN;
    output Q, QN;
endmodule
module DFKCND4 (D, CP, CN, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input D, CP, CN;
    output Q, QN;
endmodule
module DFKCNQD1 (D, CP, CN, Q);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input D, CP, CN;
    output Q;
endmodule
module DFKCNQD2 (D, CP, CN, Q);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input D, CP, CN;
    output Q;
endmodule
module DFKCNQD4 (D, CP, CN, Q);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input D, CP, CN;
    output Q;
endmodule
module DFKCSND1 (D, CP, CN, SN, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input D, CP, CN, SN;
    output Q, QN;
endmodule
module DFKCSND2 (D, CP, CN, SN, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input D, CP, CN, SN;
    output Q, QN;
endmodule
module DFKCSND4 (D, CP, CN, SN, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input D, CP, CN, SN;
    output Q, QN;
endmodule
module DFKSND1 (D, CP, SN, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input D, CP, SN;
    output Q, QN;
endmodule
module DFKSND2 (D, CP, SN, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input D, CP, SN;
    output Q, QN;
endmodule
module DFKSND4 (D, CP, SN, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input D, CP, SN;
    output Q, QN;
endmodule
module DFNCND1 (D, CPN, CDN, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input D, CPN, CDN;
    output Q, QN;
endmodule
module DFNCND2 (D, CPN, CDN, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input D, CPN, CDN;
    output Q, QN;
endmodule
module DFNCND4 (D, CPN, CDN, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input D, CPN, CDN;
    output Q, QN;
endmodule
module DFNCSND1 (D, CPN, CDN, SDN, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input D, CPN, CDN, SDN;
    output Q, QN;
endmodule
module DFNCSND2 (D, CPN, CDN, SDN, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input D, CPN, CDN, SDN;
    output Q, QN;
endmodule
module DFNCSND4 (D, CPN, CDN, SDN, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input D, CPN, CDN, SDN;
    output Q, QN;
endmodule
module DFND1 (D, CPN, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input D, CPN;
    output Q, QN;
endmodule
module DFND2 (D, CPN, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input D, CPN;
    output Q, QN;
endmodule
module DFND4 (D, CPN, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input D, CPN;
    output Q, QN;
endmodule
module DFNSND1 (D, CPN, SDN, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input D, CPN, SDN;
    output Q, QN;
endmodule
module DFNSND2 (D, CPN, SDN, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input D, CPN, SDN;
    output Q, QN;
endmodule
module DFNSND4 (D, CPN, SDN, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input D, CPN, SDN;
    output Q, QN;
endmodule
module DFQD1 (D, CP, Q);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input D, CP;
    output Q;
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
endmodule
module DFQD2 (D, CP, Q);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input D, CP;
    output Q;
endmodule
module DFQD4 (D, CP, Q);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input D, CP;
    output Q;
endmodule
module DFSND1 (D, CP, SDN, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input D, CP, SDN;
    output Q, QN;
endmodule
module DFSND2 (D, CP, SDN, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input D, CP, SDN;
    output Q, QN;
endmodule
module DFSND4 (D, CP, SDN, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input D, CP, SDN;
    output Q, QN;
endmodule
module DFSNQD1 (D, CP, SDN, Q);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input D, CP, SDN;
    output Q;
endmodule
module DFSNQD2 (D, CP, SDN, Q);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input D, CP, SDN;
    output Q;
endmodule
module DFSNQD4 (D, CP, SDN, Q);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input D, CP, SDN;
    output Q;
endmodule
module DFXD1 (DA, DB, SA, CP, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input DA, DB, SA, CP;
    output Q, QN;
endmodule
module DFXD2 (DA, DB, SA, CP, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input DA, DB, SA, CP;
    output Q, QN;
endmodule
module DFXD4 (DA, DB, SA, CP, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input DA, DB, SA, CP;
    output Q, QN;
endmodule
module DFXQD1 (DA, DB, SA, CP, Q);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input DA, DB, SA, CP;
    output Q;
endmodule
module DFXQD2 (DA, DB, SA, CP, Q);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input DA, DB, SA, CP;
    output Q;
endmodule
module DFXQD4 (DA, DB, SA, CP, Q);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input DA, DB, SA, CP;
    output Q;
endmodule
module EDFCND1 (D, E, CP, CDN, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input D, E, CP, CDN;  
    output Q, QN;
endmodule
module EDFCND2 (D, E, CP, CDN, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input D, E, CP, CDN;  
    output Q, QN;
endmodule
module EDFCND4 (D, E, CP, CDN, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input D, E, CP, CDN;  
    output Q, QN;
endmodule
module EDFCNQD1 (D, E, CP, CDN, Q);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input D, E, CP, CDN;  
    output Q;
endmodule
module EDFCNQD2 (D, E, CP, CDN, Q);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input D, E, CP, CDN;  
    output Q;
endmodule
module EDFCNQD4 (D, E, CP, CDN, Q);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input D, E, CP, CDN;  
    output Q;
endmodule
module EDFD1 (D, E, CP, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input D, E, CP;  
    output Q, QN;
endmodule
module EDFD2 (D, E, CP, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input D, E, CP;  
    output Q, QN;
endmodule
module EDFD4 (D, E, CP, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input D, E, CP;  
    output Q, QN;
endmodule
module EDFKCND1 (D, E, CP, CN, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input D, E, CP, CN;
    output Q, QN;
endmodule
module EDFKCND2 (D, E, CP, CN, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input D, E, CP, CN;
    output Q, QN;
endmodule
module EDFKCND4 (D, E, CP, CN, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input D, E, CP, CN;
    output Q, QN;
endmodule
module EDFKCNQD1 (D, E, CP, CN, Q);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input D, E, CP, CN;
    output Q;
endmodule
module EDFKCNQD2 (D, E, CP, CN, Q);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input D, E, CP, CN;
    output Q;
endmodule
module EDFKCNQD4 (D, E, CP, CN, Q);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input D, E, CP, CN;
    output Q;
endmodule
module EDFQD1 (D, E, CP, Q);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input D, E, CP;  
    output Q;
endmodule
module EDFQD2 (D, E, CP, Q);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input D, E, CP;  
    output Q;
endmodule
module EDFQD4 (D, E, CP, Q);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input D, E, CP;  
    output Q;
endmodule
module FA1D0 (A, B, CI, S, CO);
  input		A, B, CI;
  output	S, CO;
endmodule
module FA1D1 (A, B, CI, S, CO);
  input		A, B, CI;
  output	S, CO;
endmodule
module FA1D2 (A, B, CI, S, CO);
  input		A, B, CI;
  output	S, CO;
endmodule
module FA1D4 (A, B, CI, S, CO);
  input		A, B, CI;
  output	S, CO;
endmodule
module FCICIND1 (A, B, CIN, CO);
input A, B, CIN;
output CO;
endmodule
module FCICIND2 (A, B, CIN, CO);
input A, B, CIN;
output CO;
endmodule
module FCICOND1 (A, B, CI, CON);
input A, B, CI;
output CON;
endmodule
module FCICOND2 (A, B, CI, CON);
input A, B, CI;
output CON;
endmodule
module FCSICIND1 (A, B, CIN0, CIN1, CS, S, CO0, CO1);
input A, B, CIN0, CIN1, CS;
output S, CO0, CO1;
endmodule
module FCSICIND2 (A, B, CIN0, CIN1, CS, S, CO0, CO1);
input A, B, CIN0, CIN1, CS;
output S, CO0, CO1;
endmodule
module FCSICOND1 (A, B, CI0, CI1, CS, S, CON0, CON1);
input A, B, CI0, CI1, CS;
output S, CON0, CON1;
endmodule
module FCSICOND2 (A, B, CI0, CI1, CS, S, CON0, CON1);
input A, B, CI0, CI1, CS;
output S, CON0, CON1;
endmodule
module FICIND1 (A, B, CIN, S, CO);
input A, B, CIN;
output S, CO;
endmodule
module FICIND2 (A, B, CIN, S, CO);
input A, B, CIN;
output S, CO;
endmodule
module FICOND1 (A, B, CI, S, CON);
input A, B, CI;
output S, CON;
endmodule
module FICOND2 (A, B, CI, S, CON);
input A, B, CI;
output S, CON;
endmodule
module FIICOND1 (A, B, C, S, CON0, CON1);
input A, B, C;
output S, CON0, CON1;
endmodule
module FIICOND2 (A, B, C, S, CON0, CON1);
input A, B, C;
output S, CON0, CON1;
endmodule
module GAN2D1 (A1, A2, Z);
    input A1, A2;
    output Z;
endmodule
module GAN2D2 (A1, A2, Z);
    input A1, A2;
    output Z;
endmodule
module GAOI21D1 (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
endmodule
module GAOI21D2 (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
endmodule
module GAOI22D1 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
endmodule
module GBUFFD1 (I, Z);
    input I;
    output Z;
endmodule
module GBUFFD2 (I, Z);
    input I;
    output Z;
endmodule
module GBUFFD3 (I, Z);
    input I;
    output Z;
endmodule
module GBUFFD4 (I, Z);
    input I;
    output Z;
endmodule
module GBUFFD8 (I, Z);
    input I;
    output Z;
endmodule
module GDCAP;
endmodule
module GDCAP10;
endmodule
module GDCAP2;
endmodule
module GDCAP3;
endmodule
module GDCAP4;
endmodule
module GDFCNQD1 (D, CP, CDN, Q);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input D, CP, CDN;
    output Q;
endmodule
module GDFQD1 (D, CP, Q);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input D, CP;
    output Q;
endmodule
module GFILL;
endmodule
module GFILL10;
endmodule
module GFILL2;
endmodule
module GFILL3;
endmodule
module GFILL4;
endmodule
module GINVD1 (I, ZN);
    input I;
    output ZN;
endmodule
module GINVD2 (I, ZN);
    input I;
    output ZN;
endmodule
module GINVD3 (I, ZN);
    input I;
    output ZN;
endmodule
module GINVD4 (I, ZN);
    input I;
    output ZN;
endmodule
module GINVD8 (I, ZN);
    input I;
    output ZN;
endmodule
module GMUX2D1 (I0, I1, S, Z);
  input		I0, I1, S;
  output	Z;
endmodule
module GMUX2D2 (I0, I1, S, Z);
  input		I0, I1, S;
  output	Z;
endmodule
module GMUX2ND1 (I0, I1, S, ZN);
  input		 I0, I1, S;
  output	 ZN;
endmodule
module GMUX2ND2 (I0, I1, S, ZN);
  input		 I0, I1, S;
  output	 ZN;
endmodule
module GND2D1 (A1, A2, ZN);
    input A1, A2;
    output ZN;
endmodule
module GND2D2 (A1, A2, ZN);
    input A1, A2;
    output ZN;
endmodule
module GND2D3 (A1, A2, ZN);
    input A1, A2;
    output ZN;
endmodule
module GND2D4 (A1, A2, ZN);
    input A1, A2;
    output ZN;
endmodule
module GND3D1 (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
endmodule
module GND3D2 (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
endmodule
module GNR2D1 (A1, A2, ZN);
    input A1, A2;
    output ZN;
endmodule
module GNR2D2 (A1, A2, ZN);
    input A1, A2;
    output ZN;
endmodule
module GNR3D1 (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
endmodule
module GNR3D2 (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
endmodule
module GOAI21D1 (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
endmodule
module GOAI21D2 (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
endmodule
module GOR2D1 (A1, A2, Z);
    input A1, A2;
    output Z;
endmodule
module GOR2D2 (A1, A2, Z);
    input A1, A2;
    output Z;
endmodule
module GSDFCNQD1 (SI, D, SE, CP, CDN, Q);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input SI, D, SE, CP, CDN;
    output Q;
endmodule
module GTIEH (Z);
  output  Z;
endmodule
module GTIEL (ZN);
  output  ZN;
endmodule
module GXNR2D1 (A1, A2, ZN);
  input		A1, A2;
  output 	ZN;
endmodule
module GXNR2D2 (A1, A2, ZN);
  input		A1, A2;
  output 	ZN;
endmodule
module GXOR2D1 (A1, A2, Z);
  input 	A1, A2;
  output 	Z;
endmodule
module GXOR2D2 (A1, A2, Z);
  input 	A1, A2;
  output 	Z;
endmodule
module HA1D0 (A, B, S, CO);
  input	 	A, B;
  output	S, CO;
endmodule
module HA1D1 (A, B, S, CO);
  input	 	A, B;
  output	S, CO;
endmodule
module HA1D2 (A, B, S, CO);
  input	 	A, B;
  output	S, CO;
endmodule
module HA1D4 (A, B, S, CO);
  input	 	A, B;
  output	S, CO;
endmodule
module HCOSCIND1 (A, CIN, CS, S, CO);
input A, CIN, CS;
output S, CO;
endmodule
module HCOSCIND2 (A, CIN, CS, S, CO);
input A, CIN, CS;
output S, CO;
endmodule
module HCOSCOND1 (A, CI, CS, S, CON);
input A, CI, CS;
output S, CON;
endmodule
module HCOSCOND2 (A, CI, CS, S, CON);
input A, CI, CS;
output S, CON;
endmodule
module HICIND1 (A, CIN, S, CO);
input A, CIN;
output S, CO;
endmodule
module HICIND2 (A, CIN, S, CO);
input A, CIN;
output S, CO;
endmodule
module HICOND1 (A, CI, S, CON);
input A, CI;
output S, CON;
endmodule
module HICOND2 (A, CI, S, CON);
input A, CI;
output S, CON;
endmodule
module IAO21D0 (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
endmodule
module IAO21D1 (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
endmodule
module IAO21D2 (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
endmodule
module IAO21D4 (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
endmodule
module IAO22D0 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
endmodule
module IAO22D1 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
endmodule
module IAO22D2 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
endmodule
module IAO22D4 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
endmodule
module IIND4D0 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
endmodule
module IIND4D1 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
endmodule
module IIND4D2 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
endmodule
module IIND4D4 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
endmodule
module IINR4D0 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
endmodule
module IINR4D1 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
endmodule
module IINR4D2 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
endmodule
module IINR4D4 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
endmodule
module IND2D0 (A1, B1, ZN);
    input A1, B1;
    output ZN;
endmodule
module IND2D1 (A1, B1, ZN);
    input A1, B1;
    output ZN;
endmodule
module IND2D2 (A1, B1, ZN);
    input A1, B1;
    output ZN;
endmodule
module IND2D4 (A1, B1, ZN);
    input A1, B1;
    output ZN;
endmodule
module IND3D0 (A1, B1, B2, ZN);
    input A1, B1, B2;
    output ZN;
endmodule
module IND3D1 (A1, B1, B2, ZN);
    input A1, B1, B2;
    output ZN;
endmodule
module IND3D2 (A1, B1, B2, ZN);
    input A1, B1, B2;
    output ZN;
endmodule
module IND3D4 (A1, B1, B2, ZN);
    input A1, B1, B2;
    output ZN;
endmodule
module IND4D0 (A1, B1, B2, B3, ZN);
    input A1, B1, B2, B3;
    output ZN;
endmodule
module IND4D1 (A1, B1, B2, B3, ZN);
    input A1, B1, B2, B3;
    output ZN;
endmodule
module IND4D2 (A1, B1, B2, B3, ZN);
    input A1, B1, B2, B3;
    output ZN;
endmodule
module IND4D4 (A1, B1, B2, B3, ZN);
    input A1, B1, B2, B3;
    output ZN;
endmodule
module INR2D0 (A1, B1, ZN);
    input A1, B1;
    output ZN;
endmodule
module INR2D1 (A1, B1, ZN);
    input A1, B1;
    output ZN;
endmodule
module INR2D2 (A1, B1, ZN);
    input A1, B1;
    output ZN;
endmodule
module INR2D4 (A1, B1, ZN);
    input A1, B1;
    output ZN;
endmodule
module INR2XD0 (A1, B1, ZN);
    input A1, B1;
    output ZN;
endmodule
module INR2XD1 (A1, B1, ZN);
    input A1, B1;
    output ZN;
endmodule
module INR2XD2 (A1, B1, ZN);
    input A1, B1;
    output ZN;
endmodule
module INR2XD4 (A1, B1, ZN);
    input A1, B1;
    output ZN;
endmodule
module INR3D0 (A1, B1, B2, ZN);
    input A1, B1, B2;
    output ZN;
endmodule
module INR3D1 (A1, B1, B2, ZN);
    input A1, B1, B2;
    output ZN;
endmodule
module INR3D2 (A1, B1, B2, ZN);
    input A1, B1, B2;
    output ZN;
endmodule
module INR3D4 (A1, B1, B2, ZN);
    input A1, B1, B2;
    output ZN;
endmodule
module INR4D0 (A1, B1, B2, B3, ZN);
    input A1, B1, B2, B3;
    output ZN;
endmodule
module INR4D1 (A1, B1, B2, B3, ZN);
    input A1, B1, B2, B3;
    output ZN;
endmodule
module INR4D2 (A1, B1, B2, B3, ZN);
    input A1, B1, B2, B3;
    output ZN;
endmodule
module INR4D4 (A1, B1, B2, B3, ZN);
    input A1, B1, B2, B3;
    output ZN;
endmodule
module INVD0 (I, ZN);
    input I;
    output ZN;
endmodule
module INVD1 (I, ZN);
    input I;
    output ZN;
endmodule
module INVD12 (I, ZN);
    input I;
    output ZN;
endmodule
module INVD16 (I, ZN);
    input I;
    output ZN;
endmodule
module INVD2 (I, ZN);
    input I;
    output ZN;
endmodule
module INVD20 (I, ZN);
    input I;
    output ZN;
endmodule
module INVD24 (I, ZN);
    input I;
    output ZN;
endmodule
module INVD3 (I, ZN);
    input I;
    output ZN;
endmodule
module INVD4 (I, ZN);
    input I;
    output ZN;
endmodule
module INVD6 (I, ZN);
    input I;
    output ZN;
endmodule
module INVD8 (I, ZN);
    input I;
    output ZN;
endmodule
module IOA21D0 (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
endmodule
module IOA21D1 (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
endmodule
module IOA21D2 (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
endmodule
module IOA21D4 (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
endmodule
module IOA22D0 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
endmodule
module IOA22D1 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
endmodule
module IOA22D2 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
endmodule
module IOA22D4 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
endmodule
module LHCND1 (D, E, CDN, Q, QN);
    input D, E, CDN;
    output Q, QN;
endmodule
module LHCND2 (D, E, CDN, Q, QN);
    input D, E, CDN;
    output Q, QN;
endmodule
module LHCND4 (D, E, CDN, Q, QN);
    input D, E, CDN;
    output Q, QN;
endmodule
module LHCNDD1 (D, E, CDN, Q, QN);
    input D, E, CDN;
    output Q, QN;
endmodule
module LHCNDD2 (D, E, CDN, Q, QN);
    input D, E, CDN;
    output Q, QN;
endmodule
module LHCNDD4 (D, E, CDN, Q, QN);
    input D, E, CDN;
    output Q, QN;
endmodule
module LHCNDQD1 (D, E, CDN, Q);
    input D, E, CDN;
    output Q;
endmodule
module LHCNDQD2 (D, E, CDN, Q);
    input D, E, CDN;
    output Q;
endmodule
module LHCNDQD4 (D, E, CDN, Q);
    input D, E, CDN;
    output Q;
endmodule
module LHCNQD1 (D, E, CDN, Q);
    input D, E, CDN;
    output Q;
endmodule
module LHCNQD2 (D, E, CDN, Q);
    input D, E, CDN;
    output Q;
endmodule
module LHCNQD4 (D, E, CDN, Q);
    input D, E, CDN;
    output Q;
endmodule
module LHCSND1 (D, E, CDN, SDN, Q, QN);
    input D, E, CDN, SDN;
    output Q, QN;
endmodule
module LHCSND2 (D, E, CDN, SDN, Q, QN);
    input D, E, CDN, SDN;
    output Q, QN;
endmodule
module LHCSND4 (D, E, CDN, SDN, Q, QN);
    input D, E, CDN, SDN;
    output Q, QN;
endmodule
module LHCSNDD1 (D, E, CDN, SDN, Q, QN);
    input D, E, CDN, SDN;
    output Q, QN;
endmodule
module LHCSNDD2 (D, E, CDN, SDN, Q, QN);
    input D, E, CDN, SDN;
    output Q, QN;
endmodule
module LHCSNDD4 (D, E, CDN, SDN, Q, QN);
    input D, E, CDN, SDN;
    output Q, QN;
endmodule
module LHCSNDQD1 (D, E, CDN, SDN, Q);
    input D, E, CDN, SDN;
    output Q;
endmodule
module LHCSNDQD2 (D, E, CDN, SDN, Q);
    input D, E, CDN, SDN;
    output Q;
endmodule
module LHCSNDQD4 (D, E, CDN, SDN, Q);
    input D, E, CDN, SDN;
    output Q;
endmodule
module LHCSNQD1 (D, E, CDN, SDN, Q);
    input D, E, CDN, SDN;
    output Q;
endmodule
module LHCSNQD2 (D, E, CDN, SDN, Q);
    input D, E, CDN, SDN;
    output Q;
endmodule
module LHCSNQD4 (D, E, CDN, SDN, Q);
    input D, E, CDN, SDN;
    output Q;
endmodule
module LHD1 (D, E, Q, QN);
    input D, E;
    output Q, QN;
endmodule
module LHD2 (D, E, Q, QN);
    input D, E;
    output Q, QN;
endmodule
module LHD4 (D, E, Q, QN);
    input D, E;
    output Q, QN;
endmodule
module LHQD1 (D, E, Q);
    input D, E;
    output Q;
endmodule
module LHQD2 (D, E, Q);
    input D, E;
    output Q;
endmodule
module LHQD4 (D, E, Q);
    input D, E;
    output Q;
endmodule
module LHSND1 (D, E, SDN, Q, QN);
    input D, E, SDN;
    output Q, QN;
endmodule
module LHSND2 (D, E, SDN, Q, QN);
    input D, E, SDN;
    output Q, QN;
endmodule
module LHSND4 (D, E, SDN, Q, QN);
    input D, E, SDN;
    output Q, QN;
endmodule
module LHSNDD1 (D, E, SDN, Q, QN);
    input D, E, SDN;
    output Q, QN;
endmodule
module LHSNDD2 (D, E, SDN, Q, QN);
    input D, E, SDN;
    output Q, QN;
endmodule
module LHSNDD4 (D, E, SDN, Q, QN);
    input D, E, SDN;
    output Q, QN;
endmodule
module LHSNDQD1 (D, E, SDN, Q);
    input D, E, SDN;
    output Q;
endmodule
module LHSNDQD2 (D, E, SDN, Q);
    input D, E, SDN;
    output Q;
endmodule
module LHSNDQD4 (D, E, SDN, Q);
    input D, E, SDN;
    output Q;
endmodule
module LHSNQD1 (D, E, SDN, Q);
    input D, E, SDN;
    output Q;
endmodule
module LHSNQD2 (D, E, SDN, Q);
    input D, E, SDN;
    output Q;
endmodule
module LHSNQD4 (D, E, SDN, Q);
    input D, E, SDN;
    output Q;
endmodule
module LNCND1 (D, EN, CDN, Q, QN);
    input D, EN, CDN;
    output Q, QN;
endmodule
module LNCND2 (D, EN, CDN, Q, QN);
    input D, EN, CDN;
    output Q, QN;
endmodule
module LNCND4 (D, EN, CDN, Q, QN);
    input D, EN, CDN;
    output Q, QN;
endmodule
module LNCNDD1 (D, EN, CDN, Q, QN);
    input D, EN, CDN;
    output Q, QN;
endmodule
module LNCNDD2 (D, EN, CDN, Q, QN);
    input D, EN, CDN;
    output Q, QN;
endmodule
module LNCNDD4 (D, EN, CDN, Q, QN);
    input D, EN, CDN;
    output Q, QN;
endmodule
module LNCNDQD1 (D, EN, CDN, Q);
    input D, EN, CDN;
    output Q;
endmodule
module LNCNDQD2 (D, EN, CDN, Q);
    input D, EN, CDN;
    output Q;
endmodule
module LNCNDQD4 (D, EN, CDN, Q);
    input D, EN, CDN;
    output Q;
endmodule
module LNCNQD1 (D, EN, CDN, Q);
    input D, EN, CDN;
    output Q;
endmodule
module LNCNQD2 (D, EN, CDN, Q);
    input D, EN, CDN;
    output Q;
endmodule
module LNCNQD4 (D, EN, CDN, Q);
    input D, EN, CDN;
    output Q;
endmodule
module LNCSND1 (D, EN, CDN, SDN, Q, QN);
   input D, EN, CDN, SDN;
   output Q, QN;
endmodule
module LNCSND2 (D, EN, CDN, SDN, Q, QN);
   input D, EN, CDN, SDN;
   output Q, QN;
endmodule
module LNCSND4 (D, EN, CDN, SDN, Q, QN);
   input D, EN, CDN, SDN;
   output Q, QN;
endmodule
module LNCSNDD1 (D, EN, CDN, SDN, Q, QN);
   input D, EN, CDN, SDN;
   output Q, QN;
endmodule
module LNCSNDD2 (D, EN, CDN, SDN, Q, QN);
   input D, EN, CDN, SDN;
   output Q, QN;
endmodule
module LNCSNDD4 (D, EN, CDN, SDN, Q, QN);
   input D, EN, CDN, SDN;
   output Q, QN;
endmodule
module LNCSNDQD1 (D, EN, CDN, SDN, Q);
   input D, EN, CDN, SDN;
   output Q;
endmodule
module LNCSNDQD2 (D, EN, CDN, SDN, Q);
   input D, EN, CDN, SDN;
   output Q;
endmodule
module LNCSNDQD4 (D, EN, CDN, SDN, Q);
   input D, EN, CDN, SDN;
   output Q;
endmodule
module LNCSNQD1 (D, EN, CDN, SDN, Q);
   input D, EN, CDN, SDN;
   output Q;
endmodule
module LNCSNQD2 (D, EN, CDN, SDN, Q);
   input D, EN, CDN, SDN;
   output Q;
endmodule
module LNCSNQD4 (D, EN, CDN, SDN, Q);
   input D, EN, CDN, SDN;
   output Q;
endmodule
module LND1 (D, EN, Q, QN);
    input D, EN;
    output Q, QN;
endmodule
module LND2 (D, EN, Q, QN);
    input D, EN;
    output Q, QN;
endmodule
module LND4 (D, EN, Q, QN);
    input D, EN;
    output Q, QN;
endmodule
module LNQD1 (D, EN, Q);
    input D, EN;
    output Q;
endmodule
module LNQD2 (D, EN, Q);
    input D, EN;
    output Q;
endmodule
module LNQD4 (D, EN, Q);
    input D, EN;
    output Q;
endmodule
module LNSND1 (D, EN, SDN, Q, QN);
    input D, EN, SDN;
    output Q, QN;
endmodule
module LNSND2 (D, EN, SDN, Q, QN);
    input D, EN, SDN;
    output Q, QN;
endmodule
module LNSND4 (D, EN, SDN, Q, QN);
    input D, EN, SDN;
    output Q, QN;
endmodule
module LNSNDD1 (D, EN, SDN, Q, QN);
    input D, EN, SDN;
    output Q, QN;
endmodule
module LNSNDD2 (D, EN, SDN, Q, QN);
    input D, EN, SDN;
    output Q, QN;
endmodule
module LNSNDD4 (D, EN, SDN, Q, QN);
    input D, EN, SDN;
    output Q, QN;
endmodule
module LNSNDQD1 (D, EN, SDN, Q);
    input D, EN, SDN;
    output Q;
endmodule
module LNSNDQD2 (D, EN, SDN, Q);
    input D, EN, SDN;
    output Q;
endmodule
module LNSNDQD4 (D, EN, SDN, Q);
    input D, EN, SDN;
    output Q;
endmodule
module LNSNQD1 (D, EN, SDN, Q);
    input D, EN, SDN;
    output Q;
endmodule
module LNSNQD2 (D, EN, SDN, Q);
    input D, EN, SDN;
    output Q;
endmodule
module LNSNQD4 (D, EN, SDN, Q);
    input D, EN, SDN;
    output Q;
endmodule
module MAOI222D0 (A, B, C, ZN);
    input A, B, C;
    output ZN;
endmodule
module MAOI222D1 (A, B, C, ZN);
    input A, B, C;
    output ZN;
endmodule
module MAOI222D2 (A, B, C, ZN);
    input A, B, C;
    output ZN;
endmodule
module MAOI222D4 (A, B, C, ZN);
    input A, B, C;
    output ZN;
endmodule
module MAOI22D0 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
endmodule
module MAOI22D1 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
endmodule
module MAOI22D2 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
endmodule
module MAOI22D4 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
endmodule
module MOAI22D0 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
endmodule
module MOAI22D1 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
endmodule
module MOAI22D2 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
endmodule
module MOAI22D4 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
endmodule
module MUX2D0 (I0, I1, S, Z);
  input		I0, I1, S;
  output	Z;
endmodule
module MUX2D1 (I0, I1, S, Z);
  input		I0, I1, S;
  output	Z;
endmodule
module MUX2D2 (I0, I1, S, Z);
  input		I0, I1, S;
  output	Z;
endmodule
module MUX2D4 (I0, I1, S, Z);
  input		I0, I1, S;
  output	Z;
endmodule
module MUX2ND0 (I0, I1, S, ZN);
  input		 I0, I1, S;
  output	 ZN;
endmodule
module MUX2ND1 (I0, I1, S, ZN);
  input		 I0, I1, S;
  output	 ZN;
endmodule
module MUX2ND2 (I0, I1, S, ZN);
  input		 I0, I1, S;
  output	 ZN;
endmodule
module MUX2ND4 (I0, I1, S, ZN);
  input		 I0, I1, S;
  output	 ZN;
endmodule
module MUX3D0 (I0, I1, I2, S0, S1, Z);
  input		I0, I1, I2, S0, S1;
  output	Z;
endmodule
module MUX3D1 (I0, I1, I2, S0, S1, Z);
  input		I0, I1, I2, S0, S1;
  output	Z;
endmodule
module MUX3D2 (I0, I1, I2, S0, S1, Z);
  input		I0, I1, I2, S0, S1;
  output	Z;
endmodule
module MUX3D4 (I0, I1, I2, S0, S1, Z);
  input		I0, I1, I2, S0, S1;
  output	Z;
endmodule
module MUX3ND0 (I0, I1, I2, S0, S1, ZN);
  input 	I0, I1, I2, S0, S1;
  output 	ZN;
endmodule
module MUX3ND1 (I0, I1, I2, S0, S1, ZN);
  input 	I0, I1, I2, S0, S1;
  output 	ZN;
endmodule
module MUX3ND2 (I0, I1, I2, S0, S1, ZN);
  input 	I0, I1, I2, S0, S1;
  output 	ZN;
endmodule
module MUX3ND4 (I0, I1, I2, S0, S1, ZN);
  input 	I0, I1, I2, S0, S1;
  output 	ZN;
endmodule
module MUX4D0 (I0, I1, I2, I3, S0, S1, Z);
  input		 I0, I1, I2, I3, S0, S1;
  output	 Z;
endmodule
module MUX4D1 (I0, I1, I2, I3, S0, S1, Z);
  input		 I0, I1, I2, I3, S0, S1;
  output	 Z;
endmodule
module MUX4D2 (I0, I1, I2, I3, S0, S1, Z);
  input		 I0, I1, I2, I3, S0, S1;
  output	 Z;
endmodule
module MUX4D4 (I0, I1, I2, I3, S0, S1, Z);
  input		 I0, I1, I2, I3, S0, S1;
  output	 Z;
endmodule
module MUX4ND0 (I0, I1, I2, I3, S0, S1, ZN);
  input		 I0, I1, I2, I3, S0, S1;
  output	 ZN;
endmodule
module MUX4ND1 (I0, I1, I2, I3, S0, S1, ZN);
  input		 I0, I1, I2, I3, S0, S1;
  output	 ZN;
endmodule
module MUX4ND2 (I0, I1, I2, I3, S0, S1, ZN);
  input		 I0, I1, I2, I3, S0, S1;
  output	 ZN;
endmodule
module MUX4ND4 (I0, I1, I2, I3, S0, S1, ZN);
  input		 I0, I1, I2, I3, S0, S1;
  output	 ZN;
endmodule
module ND2D0 (A1, A2, ZN);
    input A1, A2;
    output ZN;
endmodule
module ND2D1 (A1, A2, ZN);
    input A1, A2;
    output ZN;
endmodule
module ND2D2 (A1, A2, ZN);
    input A1, A2;
    output ZN;
endmodule
module ND2D3 (A1, A2, ZN);
    input A1, A2;
    output ZN;
endmodule
module ND2D4 (A1, A2, ZN);
    input A1, A2;
    output ZN;
endmodule
module ND2D8 (A1, A2, ZN);
    input A1, A2;
    output ZN;
endmodule
module ND3D0 (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
endmodule
module ND3D1 (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
endmodule
module ND3D2 (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
endmodule
module ND3D3 (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
endmodule
module ND3D4 (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
endmodule
module ND3D8 (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
endmodule
module ND4D0 (A1, A2, A3, A4, ZN);
    input A1, A2, A3, A4;
    output ZN;
endmodule
module ND4D1 (A1, A2, A3, A4, ZN);
    input A1, A2, A3, A4;
    output ZN;
endmodule
module ND4D2 (A1, A2, A3, A4, ZN);
    input A1, A2, A3, A4;
    output ZN;
endmodule
module ND4D3 (A1, A2, A3, A4, ZN);
    input A1, A2, A3, A4;
    output ZN;
endmodule
module ND4D4 (A1, A2, A3, A4, ZN);
    input A1, A2, A3, A4;
    output ZN;
endmodule
module ND4D8 (A1, A2, A3, A4, ZN);
    input A1, A2, A3, A4;
    output ZN;
endmodule
module NR2D0 (A1, A2, ZN);
    input A1, A2;
    output ZN;
endmodule
module NR2D1 (A1, A2, ZN);
    input A1, A2;
    output ZN;
endmodule
module NR2D2 (A1, A2, ZN);
    input A1, A2;
    output ZN;
endmodule
module NR2D3 (A1, A2, ZN);
    input A1, A2;
    output ZN;
endmodule
module NR2D4 (A1, A2, ZN);
    input A1, A2;
    output ZN;
endmodule
module NR2D8 (A1, A2, ZN);
    input A1, A2;
    output ZN;
endmodule
module NR2XD0 (A1, A2, ZN);
    input A1, A2;
    output ZN;
endmodule
module NR2XD1 (A1, A2, ZN);
    input A1, A2;
    output ZN;
endmodule
module NR2XD2 (A1, A2, ZN);
    input A1, A2;
    output ZN;
endmodule
module NR2XD3 (A1, A2, ZN);
    input A1, A2;
    output ZN;
endmodule
module NR2XD4 (A1, A2, ZN);
    input A1, A2;
    output ZN;
endmodule
module NR2XD8 (A1, A2, ZN);
    input A1, A2;
    output ZN;
endmodule
module NR3D0 (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
endmodule
module NR3D1 (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
endmodule
module NR3D2 (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
endmodule
module NR3D3 (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
endmodule
module NR3D4 (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
endmodule
module NR3D8 (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
endmodule
module NR4D0 (A1, A2, A3, A4, ZN);
    input A1, A2, A3, A4;
    output ZN;
endmodule
module NR4D1 (A1, A2, A3, A4, ZN);
    input A1, A2, A3, A4;
    output ZN;
endmodule
module NR4D2 (A1, A2, A3, A4, ZN);
    input A1, A2, A3, A4;
    output ZN;
endmodule
module NR4D3 (A1, A2, A3, A4, ZN);
    input A1, A2, A3, A4;
    output ZN;
endmodule
module NR4D4 (A1, A2, A3, A4, ZN);
    input A1, A2, A3, A4;
    output ZN;
endmodule
module NR4D8 (A1, A2, A3, A4, ZN);
    input A1, A2, A3, A4;
    output ZN;
endmodule
module OA211D0 (A1, A2, B, C, Z);
    input A1, A2, B, C;
    output Z;
endmodule
module OA211D1 (A1, A2, B, C, Z);
    input A1, A2, B, C;
    output Z;
endmodule
module OA211D2 (A1, A2, B, C, Z);
    input A1, A2, B, C;
    output Z;
endmodule
module OA211D4 (A1, A2, B, C, Z);
    input A1, A2, B, C;
    output Z;
endmodule
module OA21D0 (A1, A2, B, Z);
    input A1, A2, B;
    output Z;
endmodule
module OA21D1 (A1, A2, B, Z);
    input A1, A2, B;
    output Z;
endmodule
module OA21D2 (A1, A2, B, Z);
    input A1, A2, B;
    output Z;
endmodule
module OA21D4 (A1, A2, B, Z);
    input A1, A2, B;
    output Z;
endmodule
module OA221D0 (A1, A2, B1, B2, C, Z);
    input A1, A2, B1, B2, C;
    output Z;
endmodule
module OA221D1 (A1, A2, B1, B2, C, Z);
    input A1, A2, B1, B2, C;
    output Z;
endmodule
module OA221D2 (A1, A2, B1, B2, C, Z);
    input A1, A2, B1, B2, C;
    output Z;
endmodule
module OA221D4 (A1, A2, B1, B2, C, Z);
    input A1, A2, B1, B2, C;
    output Z;
endmodule
module OA222D0 (A1, A2, B1, B2, C1, C2, Z);
    input A1, A2, B1, B2, C1, C2;
    output Z;
endmodule
module OA222D1 (A1, A2, B1, B2, C1, C2, Z);
    input A1, A2, B1, B2, C1, C2;
    output Z;
endmodule
module OA222D2 (A1, A2, B1, B2, C1, C2, Z);
    input A1, A2, B1, B2, C1, C2;
    output Z;
endmodule
module OA222D4 (A1, A2, B1, B2, C1, C2, Z);
    input A1, A2, B1, B2, C1, C2;
    output Z;
endmodule
module OA22D0 (A1, A2, B1, B2, Z);
    input A1, A2, B1, B2;
    output Z;
endmodule
module OA22D1 (A1, A2, B1, B2, Z);
    input A1, A2, B1, B2;
    output Z;
endmodule
module OA22D2 (A1, A2, B1, B2, Z);
    input A1, A2, B1, B2;
    output Z;
endmodule
module OA22D4 (A1, A2, B1, B2, Z);
    input A1, A2, B1, B2;
    output Z;
endmodule
module OA31D0 (A1, A2, A3, B, Z);
    input A1, A2, A3, B;
    output Z;
endmodule
module OA31D1 (A1, A2, A3, B, Z);
    input A1, A2, A3, B;
    output Z;
endmodule
module OA31D2 (A1, A2, A3, B, Z);
    input A1, A2, A3, B;
    output Z;
endmodule
module OA31D4 (A1, A2, A3, B, Z);
    input A1, A2, A3, B;
    output Z;
endmodule
module OA32D0 (A1, A2, A3, B1, B2, Z);
    input A1, A2, A3, B1, B2;
    output Z;
endmodule
module OA32D1 (A1, A2, A3, B1, B2, Z);
    input A1, A2, A3, B1, B2;
    output Z;
endmodule
module OA32D2 (A1, A2, A3, B1, B2, Z);
    input A1, A2, A3, B1, B2;
    output Z;
endmodule
module OA32D4 (A1, A2, A3, B1, B2, Z);
    input A1, A2, A3, B1, B2;
    output Z;
endmodule
module OA33D0 (A1, A2, A3, B1, B2, B3, Z);
    input A1, A2, A3, B1, B2, B3;
    output Z;
endmodule
module OA33D1 (A1, A2, A3, B1, B2, B3, Z);
    input A1, A2, A3, B1, B2, B3;
    output Z;
endmodule
module OA33D2 (A1, A2, A3, B1, B2, B3, Z);
    input A1, A2, A3, B1, B2, B3;
    output Z;
endmodule
module OA33D4 (A1, A2, A3, B1, B2, B3, Z);
    input A1, A2, A3, B1, B2, B3;
    output Z;
endmodule
module OAI211D0 (A1, A2, B, C, ZN);
    input A1, A2, B, C;
    output ZN;
endmodule
module OAI211D1 (A1, A2, B, C, ZN);
    input A1, A2, B, C;
    output ZN;
endmodule
module OAI211D2 (A1, A2, B, C, ZN);
    input A1, A2, B, C;
    output ZN;
endmodule
module OAI211D4 (A1, A2, B, C, ZN);
    input A1, A2, B, C;
    output ZN;
endmodule
module OAI21D0 (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
endmodule
module OAI21D1 (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
endmodule
module OAI21D2 (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
endmodule
module OAI21D4 (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
endmodule
module OAI221D0 (A1, A2, B1, B2, C, ZN);
    input A1, A2, B1, B2, C;
    output ZN;
endmodule
module OAI221D1 (A1, A2, B1, B2, C, ZN);
    input A1, A2, B1, B2, C;
    output ZN;
endmodule
module OAI221D2 (A1, A2, B1, B2, C, ZN);
    input A1, A2, B1, B2, C;
    output ZN;
endmodule
module OAI221D4 (A1, A2, B1, B2, C, ZN);
    input A1, A2, B1, B2, C;
    output ZN;
endmodule
module OAI221XD4 (A1, A2, B1, B2, C, ZN);
    input A1, A2, B1, B2, C;
    output ZN;
endmodule
module OAI222D0 (A1, A2, B1, B2, C1, C2, ZN);
    input A1, A2, B1, B2, C1, C2;
    output ZN;
endmodule
module OAI222D1 (A1, A2, B1, B2, C1, C2, ZN);
    input A1, A2, B1, B2, C1, C2;
    output ZN;
endmodule
module OAI222D2 (A1, A2, B1, B2, C1, C2, ZN);
    input A1, A2, B1, B2, C1, C2;
    output ZN;
endmodule
module OAI222D4 (A1, A2, B1, B2, C1, C2, ZN);
    input A1, A2, B1, B2, C1, C2;
    output ZN;
endmodule
module OAI222XD4 (A1, A2, B1, B2, C1, C2, ZN);
    input A1, A2, B1, B2, C1, C2;
    output ZN;
endmodule
module OAI22D0 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
endmodule
module OAI22D1 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
endmodule
module OAI22D2 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
endmodule
module OAI22D4 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
endmodule
module OAI31D0 (A1, A2, A3, B, ZN);
    input A1, A2, A3, B;
    output ZN;
endmodule
module OAI31D1 (A1, A2, A3, B, ZN);
    input A1, A2, A3, B;
    output ZN;
endmodule
module OAI31D2 (A1, A2, A3, B, ZN);
    input A1, A2, A3, B;
    output ZN;
endmodule
module OAI31D4 (A1, A2, A3, B, ZN);
    input A1, A2, A3, B;
    output ZN;
endmodule
module OAI32D0 (A1, A2, A3, B1, B2, ZN);
    input A1, A2, A3, B1, B2;
    output ZN;
endmodule
module OAI32D1 (A1, A2, A3, B1, B2, ZN);
    input A1, A2, A3, B1, B2;
    output ZN;
endmodule
module OAI32D2 (A1, A2, A3, B1, B2, ZN);
    input A1, A2, A3, B1, B2;
    output ZN;
endmodule
module OAI32D4 (A1, A2, A3, B1, B2, ZN);
    input A1, A2, A3, B1, B2;
    output ZN;
endmodule
module OAI32XD4 (A1, A2, A3, B1, B2, ZN);
    input A1, A2, A3, B1, B2;
    output ZN;
endmodule
module OAI33D0 (A1, A2, A3, B1, B2, B3, ZN);
    input A1, A2, A3, B1, B2, B3;
    output ZN;
endmodule
module OAI33D1 (A1, A2, A3, B1, B2, B3, ZN);
    input A1, A2, A3, B1, B2, B3;
    output ZN;
endmodule
module OAI33D2 (A1, A2, A3, B1, B2, B3, ZN);
    input A1, A2, A3, B1, B2, B3;
    output ZN;
endmodule
module OAI33D4 (A1, A2, A3, B1, B2, B3, ZN);
    input A1, A2, A3, B1, B2, B3;
    output ZN;
endmodule
module OAI33XD4 (A1, A2, A3, B1, B2, B3, ZN);
    input A1, A2, A3, B1, B2, B3;
    output ZN;
endmodule
module OD25DCAP16;
endmodule
module OD25DCAP32;
endmodule
module OD25DCAP64;
endmodule
module OR2D0 (A1, A2, Z);
    input A1, A2;
    output Z;
endmodule
module OR2D1 (A1, A2, Z);
    input A1, A2;
    output Z;
endmodule
module OR2D2 (A1, A2, Z);
    input A1, A2;
    output Z;
endmodule
module OR2D4 (A1, A2, Z);
    input A1, A2;
    output Z;
endmodule
module OR2D8 (A1, A2, Z);
    input A1, A2;
    output Z;
endmodule
module OR2XD1 (A1, A2, Z);
    input A1, A2;
    output Z;
endmodule
module OR3D0 (A1, A2, A3, Z);
    input A1, A2, A3;
    output Z;
endmodule
module OR3D1 (A1, A2, A3, Z);
    input A1, A2, A3;
    output Z;
endmodule
module OR3D2 (A1, A2, A3, Z);
    input A1, A2, A3;
    output Z;
endmodule
module OR3D4 (A1, A2, A3, Z);
    input A1, A2, A3;
    output Z;
endmodule
module OR3D8 (A1, A2, A3, Z);
    input A1, A2, A3;
    output Z;
endmodule
module OR3XD1 (A1, A2, A3, Z);
    input A1, A2, A3;
    output Z;
endmodule
module OR4D0 (A1, A2, A3, A4, Z);
    input A1, A2, A3, A4;
    output Z;
endmodule
module OR4D1 (A1, A2, A3, A4, Z);
    input A1, A2, A3, A4;
    output Z;
endmodule
module OR4D2 (A1, A2, A3, A4, Z);
    input A1, A2, A3, A4;
    output Z;
endmodule
module OR4D4 (A1, A2, A3, A4, Z);
    input A1, A2, A3, A4;
    output Z;
endmodule
module OR4D8 (A1, A2, A3, A4, Z);
    input A1, A2, A3, A4;
    output Z;
endmodule
module OR4XD1 (A1, A2, A3, A4, Z);
    input A1, A2, A3, A4;
    output Z;
endmodule
module SDFCND0 (SI, D, SE, CP, CDN, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input SI, D, SE, CP, CDN;
    output Q, QN;
endmodule
module SDFCND1 (SI, D, SE, CP, CDN, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input SI, D, SE, CP, CDN;
    output Q, QN;
endmodule
module SDFCND2 (SI, D, SE, CP, CDN, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input SI, D, SE, CP, CDN;
    output Q, QN;
endmodule
module SDFCND4 (SI, D, SE, CP, CDN, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input SI, D, SE, CP, CDN;
    output Q, QN;
endmodule
module SDFCNQD0 (SI, D, SE, CP, CDN, Q);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input SI, D, SE, CP, CDN;
    output Q;
endmodule
module SDFCNQD1 (SI, D, SE, CP, CDN, Q);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input SI, D, SE, CP, CDN;
    output Q;
endmodule
module SDFCNQD2 (SI, D, SE, CP, CDN, Q);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input SI, D, SE, CP, CDN;
    output Q;
endmodule
module SDFCNQD4 (SI, D, SE, CP, CDN, Q);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input SI, D, SE, CP, CDN;
    output Q;
endmodule
module SDFCSND0 (SI, D, SE, CP, CDN, SDN, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input SI, D, SE, CP, CDN, SDN;
    output Q, QN;
endmodule
module SDFCSND1 (SI, D, SE, CP, CDN, SDN, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input SI, D, SE, CP, CDN, SDN;
    output Q, QN;
endmodule
module SDFCSND2 (SI, D, SE, CP, CDN, SDN, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input SI, D, SE, CP, CDN, SDN;
    output Q, QN;
endmodule
module SDFCSND4 (SI, D, SE, CP, CDN, SDN, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input SI, D, SE, CP, CDN, SDN;
    output Q, QN;
endmodule
module SDFCSNQD0 (SI, D, SE, CP, CDN, SDN, Q);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input SI, D, SE, CP, CDN, SDN;
    output Q;
endmodule
module SDFCSNQD1 (SI, D, SE, CP, CDN, SDN, Q);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input SI, D, SE, CP, CDN, SDN;
    output Q;
endmodule
module SDFCSNQD2 (SI, D, SE, CP, CDN, SDN, Q);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input SI, D, SE, CP, CDN, SDN;
    output Q;
endmodule
module SDFCSNQD4 (SI, D, SE, CP, CDN, SDN, Q);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input SI, D, SE, CP, CDN, SDN;
    output Q;
endmodule
module SDFD0 (SI, D, SE, CP, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input SI, D, SE, CP;
    output Q, QN;
endmodule
module SDFD1 (SI, D, SE, CP, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input SI, D, SE, CP;
    output Q, QN;
endmodule
module SDFD2 (SI, D, SE, CP, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input SI, D, SE, CP;
    output Q, QN;
endmodule
module SDFD4 (SI, D, SE, CP, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input SI, D, SE, CP;
    output Q, QN;
endmodule
module SDFKCND0 (SI, D, SE, CP, CN, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input SI, D, SE, CP, CN;
    output Q, QN;
endmodule
module SDFKCND1 (SI, D, SE, CP, CN, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input SI, D, SE, CP, CN;
    output Q, QN;
endmodule
module SDFKCND2 (SI, D, SE, CP, CN, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input SI, D, SE, CP, CN;
    output Q, QN;
endmodule
module SDFKCND4 (SI, D, SE, CP, CN, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input SI, D, SE, CP, CN;
    output Q, QN;
endmodule
module SDFKCNQD0 (SI, D, SE, CP, CN, Q);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input SI, D, SE, CP, CN;
    output Q;
endmodule
module SDFKCNQD1 (SI, D, SE, CP, CN, Q);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input SI, D, SE, CP, CN;
    output Q;
endmodule
module SDFKCNQD2 (SI, D, SE, CP, CN, Q);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input SI, D, SE, CP, CN;
    output Q;
endmodule
module SDFKCNQD4 (SI, D, SE, CP, CN, Q);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input SI, D, SE, CP, CN;
    output Q;
endmodule
module SDFKCSND0 (SI, D, SE, CP, CN, SN, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input SI, D, SE, CP, CN, SN;
    output Q, QN;
endmodule
module SDFKCSND1 (SI, D, SE, CP, CN, SN, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input SI, D, SE, CP, CN, SN;
    output Q, QN;
endmodule
module SDFKCSND2 (SI, D, SE, CP, CN, SN, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input SI, D, SE, CP, CN, SN;
    output Q, QN;
endmodule
module SDFKCSND4 (SI, D, SE, CP, CN, SN, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input SI, D, SE, CP, CN, SN;
    output Q, QN;
endmodule
module SDFKCSNQD0 (SI, D, SE, CP, CN, SN, Q);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input SI, D, SE, CP, CN, SN;
    output Q;
endmodule
module SDFKCSNQD1 (SI, D, SE, CP, CN, SN, Q);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input SI, D, SE, CP, CN, SN;
    output Q;
endmodule
module SDFKCSNQD2 (SI, D, SE, CP, CN, SN, Q);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input SI, D, SE, CP, CN, SN;
    output Q;
endmodule
module SDFKCSNQD4 (SI, D, SE, CP, CN, SN, Q);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input SI, D, SE, CP, CN, SN;
    output Q;
endmodule
module SDFKSND0 (SI, D, SE, CP, SN, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input SI, D, SE, CP, SN;
    output Q, QN;
endmodule
module SDFKSND1 (SI, D, SE, CP, SN, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input SI, D, SE, CP, SN;
    output Q, QN;
endmodule
module SDFKSND2 (SI, D, SE, CP, SN, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input SI, D, SE, CP, SN;
    output Q, QN;
endmodule
module SDFKSND4 (SI, D, SE, CP, SN, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input SI, D, SE, CP, SN;
    output Q, QN;
endmodule
module SDFKSNQD0 (SI, D, SE, CP, SN, Q);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input SI, D, SE, CP, SN;
    output Q;
endmodule
module SDFKSNQD1 (SI, D, SE, CP, SN, Q);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input SI, D, SE, CP, SN;
    output Q;
endmodule
module SDFKSNQD2 (SI, D, SE, CP, SN, Q);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input SI, D, SE, CP, SN;
    output Q;
endmodule
module SDFKSNQD4 (SI, D, SE, CP, SN, Q);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input SI, D, SE, CP, SN;
    output Q;
endmodule
module SDFNCND0 (SI, D, SE, CPN, CDN, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input SI, D, SE, CPN, CDN;
    output Q, QN;
endmodule
module SDFNCND1 (SI, D, SE, CPN, CDN, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input SI, D, SE, CPN, CDN;
    output Q, QN;
endmodule
module SDFNCND2 (SI, D, SE, CPN, CDN, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input SI, D, SE, CPN, CDN;
    output Q, QN;
endmodule
module SDFNCND4 (SI, D, SE, CPN, CDN, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input SI, D, SE, CPN, CDN;
    output Q, QN;
endmodule
module SDFNCSND0 (SI, D, SE, CPN, CDN, SDN, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input SI, D, SE, CPN, CDN, SDN;
    output Q, QN;
endmodule
module SDFNCSND1 (SI, D, SE, CPN, CDN, SDN, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input SI, D, SE, CPN, CDN, SDN;
    output Q, QN;
endmodule
module SDFNCSND2 (SI, D, SE, CPN, CDN, SDN, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input SI, D, SE, CPN, CDN, SDN;
    output Q, QN;
endmodule
module SDFNCSND4 (SI, D, SE, CPN, CDN, SDN, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input SI, D, SE, CPN, CDN, SDN;
    output Q, QN;
endmodule
module SDFND0 (SI, D, SE, CPN, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input SI, D, SE, CPN;
    output Q, QN;
endmodule
module SDFND1 (SI, D, SE, CPN, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input SI, D, SE, CPN;
    output Q, QN;
endmodule
module SDFND2 (SI, D, SE, CPN, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input SI, D, SE, CPN;
    output Q, QN;
endmodule
module SDFND4 (SI, D, SE, CPN, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input SI, D, SE, CPN;
    output Q, QN;
endmodule
module SDFNSND0 (SI, D, SE, CPN, SDN, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input SI, D, SE, CPN, SDN;
    output Q, QN;
endmodule
module SDFNSND1 (SI, D, SE, CPN, SDN, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input SI, D, SE, CPN, SDN;
    output Q, QN;
endmodule
module SDFNSND2 (SI, D, SE, CPN, SDN, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input SI, D, SE, CPN, SDN;
    output Q, QN;
endmodule
module SDFNSND4 (SI, D, SE, CPN, SDN, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input SI, D, SE, CPN, SDN;
    output Q, QN;
endmodule
module SDFQD0 (SI, D, SE, CP, Q);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input SI, D, SE, CP;
    output Q;
endmodule
module SDFQD1 (SI, D, SE, CP, Q);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input SI, D, SE, CP;
    output Q;
endmodule
module SDFQD2 (SI, D, SE, CP, Q);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input SI, D, SE, CP;
    output Q;
endmodule
module SDFQD4 (SI, D, SE, CP, Q);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input SI, D, SE, CP;
    output Q;
endmodule
module SDFQND0 (SI, D, SE, CP, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input SI, D, SE, CP;
    output QN;
endmodule
module SDFQND1 (SI, D, SE, CP, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input SI, D, SE, CP;
    output QN;
endmodule
module SDFQND2 (SI, D, SE, CP, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input SI, D, SE, CP;
    output QN;
endmodule
module SDFQND4 (SI, D, SE, CP, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input SI, D, SE, CP;
    output QN;
endmodule
module SDFSND0 (SI, D, SE, CP, SDN, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input SI, D, SE, CP, SDN;
    output Q, QN;
endmodule
module SDFSND1 (SI, D, SE, CP, SDN, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input SI, D, SE, CP, SDN;
    output Q, QN;
endmodule
module SDFSND2 (SI, D, SE, CP, SDN, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input SI, D, SE, CP, SDN;
    output Q, QN;
endmodule
module SDFSND4 (SI, D, SE, CP, SDN, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input SI, D, SE, CP, SDN;
    output Q, QN;
endmodule
module SDFSNQD0 (SI, D, SE, CP, SDN, Q);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input SI, D, SE, CP, SDN;
    output Q;
endmodule
module SDFSNQD1 (SI, D, SE, CP, SDN, Q);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input SI, D, SE, CP, SDN;
    output Q;
endmodule
module SDFSNQD2 (SI, D, SE, CP, SDN, Q);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input SI, D, SE, CP, SDN;
    output Q;
endmodule
module SDFSNQD4 (SI, D, SE, CP, SDN, Q);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input SI, D, SE, CP, SDN;
    output Q;
endmodule
module SDFXD0 (DA, DB, SA, SI, SE, CP, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input DA, DB, SA, SI, SE, CP;
    output Q, QN;
endmodule
module SDFXD1 (DA, DB, SA, SI, SE, CP, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input DA, DB, SA, SI, SE, CP;
    output Q, QN;
endmodule
module SDFXD2 (DA, DB, SA, SI, SE, CP, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input DA, DB, SA, SI, SE, CP;
    output Q, QN;
endmodule
module SDFXD4 (DA, DB, SA, SI, SE, CP, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input DA, DB, SA, SI, SE, CP;
    output Q, QN;
endmodule
module SDFXQD0 (DA, DB, SA, SI, SE, CP, Q);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input DA, DB, SA, SI, SE, CP;
    output Q;
endmodule
module SDFXQD1 (DA, DB, SA, SI, SE, CP, Q);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input DA, DB, SA, SI, SE, CP;
    output Q;
endmodule
module SDFXQD2 (DA, DB, SA, SI, SE, CP, Q);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input DA, DB, SA, SI, SE, CP;
    output Q;
endmodule
module SDFXQD4 (DA, DB, SA, SI, SE, CP, Q);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input DA, DB, SA, SI, SE, CP;
    output Q;
endmodule
module SEDFCND0 (E, SE, CP, SI, D, CDN, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input E, SE, CP, SI, D, CDN; 
    output Q, QN;
endmodule
module SEDFCND1 (E, SE, CP, SI, D, CDN, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input E, SE, CP, SI, D, CDN; 
    output Q, QN;
endmodule
module SEDFCND2 (E, SE, CP, SI, D, CDN, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input E, SE, CP, SI, D, CDN; 
    output Q, QN;
endmodule
module SEDFCND4 (E, SE, CP, SI, D, CDN, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input E, SE, CP, SI, D, CDN; 
    output Q, QN;
endmodule
module SEDFCNQD0 (E, SE, CP, SI, D, CDN, Q);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input E, SE, CP, SI, D, CDN; 
    output Q;
endmodule
module SEDFCNQD1 (E, SE, CP, SI, D, CDN, Q);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input E, SE, CP, SI, D, CDN; 
    output Q;
endmodule
module SEDFCNQD2 (E, SE, CP, SI, D, CDN, Q);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input E, SE, CP, SI, D, CDN; 
    output Q;
endmodule
module SEDFCNQD4 (E, SE, CP, SI, D, CDN, Q);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input E, SE, CP, SI, D, CDN; 
    output Q;
endmodule
module SEDFD0 (E, SE, CP, SI, D, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input E, SE, CP, SI, D; 
    output Q, QN;
endmodule
module SEDFD1 (E, SE, CP, SI, D, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input E, SE, CP, SI, D; 
    output Q, QN;
endmodule
module SEDFD2 (E, SE, CP, SI, D, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input E, SE, CP, SI, D; 
    output Q, QN;
endmodule
module SEDFD4 (E, SE, CP, SI, D, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input E, SE, CP, SI, D; 
    output Q, QN;
endmodule
module SEDFKCND0 (SI, D, E, SE, CP, CN, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input SI, D, SE, CP, CN, E;
    output Q, QN;
endmodule
module SEDFKCND1 (SI, D, E, SE, CP, CN, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input SI, D, SE, CP, CN, E;
    output Q, QN;
endmodule
module SEDFKCND2 (SI, D, E, SE, CP, CN, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input SI, D, SE, CP, CN, E;
    output Q, QN;
endmodule
module SEDFKCND4 (SI, D, E, SE, CP, CN, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input SI, D, SE, CP, CN, E;
    output Q, QN;
endmodule
module SEDFKCNQD0 (SI, D, E, SE, CP, CN, Q);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input SI, D, SE, CP, CN, E;
    output Q;
endmodule
module SEDFKCNQD1 (SI, D, E, SE, CP, CN, Q);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input SI, D, SE, CP, CN, E;
    output Q;
endmodule
module SEDFKCNQD2 (SI, D, E, SE, CP, CN, Q);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input SI, D, SE, CP, CN, E;
    output Q;
endmodule
module SEDFKCNQD4 (SI, D, E, SE, CP, CN, Q);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input SI, D, SE, CP, CN, E;
    output Q;
endmodule
module SEDFQD0 (E, SE, CP, SI, D, Q);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input E, SE, CP, SI, D; 
    output Q;
endmodule
module SEDFQD1 (E, SE, CP, SI, D, Q);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input E, SE, CP, SI, D; 
    output Q;
endmodule
module SEDFQD2 (E, SE, CP, SI, D, Q);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input E, SE, CP, SI, D; 
    output Q;
endmodule
module SEDFQD4 (E, SE, CP, SI, D, Q);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input E, SE, CP, SI, D; 
    output Q;
endmodule
module SEDFQND0 (E, SE, CP, SI, D, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input E, SE, CP, SI, D; 
    output QN;
endmodule
module SEDFQND1 (E, SE, CP, SI, D, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input E, SE, CP, SI, D; 
    output QN;
endmodule
module SEDFQND2 (E, SE, CP, SI, D, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input E, SE, CP, SI, D; 
    output QN;
endmodule
module SEDFQND4 (E, SE, CP, SI, D, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input E, SE, CP, SI, D; 
    output QN;
endmodule
module SEDFQNXD0 (E, SE, CP, SI, D, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input E, SE, CP, SI, D; 
    output QN;
endmodule
module SEDFQNXD1 (E, SE, CP, SI, D, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input E, SE, CP, SI, D; 
    output QN;
endmodule
module SEDFQNXD2 (E, SE, CP, SI, D, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input E, SE, CP, SI, D; 
    output QN;
endmodule
module SEDFQNXD4 (E, SE, CP, SI, D, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input E, SE, CP, SI, D; 
    output QN;
endmodule
module SEDFQXD0 (E, SE, CP, SI, D, Q);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input E, SE, CP, SI, D; 
    output Q;
endmodule
module SEDFQXD1 (E, SE, CP, SI, D, Q);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input E, SE, CP, SI, D; 
    output Q;
endmodule
module SEDFQXD2 (E, SE, CP, SI, D, Q);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input E, SE, CP, SI, D; 
    output Q;
endmodule
module SEDFQXD4 (E, SE, CP, SI, D, Q);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input E, SE, CP, SI, D; 
    output Q;
endmodule
module SEDFXD0 (E, SE, CP, SI, D, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input E, SE, CP, SI, D; 
    output Q, QN;
endmodule
module SEDFXD1 (E, SE, CP, SI, D, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input E, SE, CP, SI, D; 
    output Q, QN;
endmodule
module SEDFXD2 (E, SE, CP, SI, D, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input E, SE, CP, SI, D; 
    output Q, QN;
endmodule
module SEDFXD4 (E, SE, CP, SI, D, Q, QN);
    // tmrg seu_reset CDN
    // tmrg seu_set   SDN
    input E, SE, CP, SI, D; 
    output Q, QN;
endmodule
module TIEH (Z);
  output  Z;
endmodule
module TIEL (ZN);
  output  ZN;
endmodule
module XNR2D0 (A1, A2, ZN);
  input		A1, A2;
  output 	ZN;
endmodule
module XNR2D1 (A1, A2, ZN);
  input		A1, A2;
  output 	ZN;
endmodule
module XNR2D2 (A1, A2, ZN);
  input		A1, A2;
  output 	ZN;
endmodule
module XNR2D4 (A1, A2, ZN);
  input		A1, A2;
  output 	ZN;
endmodule
module XNR3D0 (A1, A2, A3, ZN);
  input A1, A2, A3;
  output ZN;
endmodule
module XNR3D1 (A1, A2, A3, ZN);
  input A1, A2, A3;
  output ZN;
endmodule
module XNR3D2 (A1, A2, A3, ZN);
  input A1, A2, A3;
  output ZN;
endmodule
module XNR3D4 (A1, A2, A3, ZN);
  input A1, A2, A3;
  output ZN;
endmodule
module XNR4D0 (A1, A2, A3, A4, ZN);
  input 	A1, A2, A3, A4;
  output 	ZN;
endmodule
module XNR4D1 (A1, A2, A3, A4, ZN);
  input 	A1, A2, A3, A4;
  output 	ZN;
endmodule
module XNR4D2 (A1, A2, A3, A4, ZN);
  input 	A1, A2, A3, A4;
  output 	ZN;
endmodule
module XNR4D4 (A1, A2, A3, A4, ZN);
  input 	A1, A2, A3, A4;
  output 	ZN;
endmodule
module XOR2D0 (A1, A2, Z);
  input 	A1, A2;
  output 	Z;
endmodule
module XOR2D1 (A1, A2, Z);
  input 	A1, A2;
  output 	Z;
endmodule
module XOR2D2 (A1, A2, Z);
  input 	A1, A2;
  output 	Z;
endmodule
module XOR2D4 (A1, A2, Z);
  input 	A1, A2;
  output 	Z;
endmodule
module XOR3D0 (A1, A2, A3, Z);
  input A1, A2, A3;
  output Z;
endmodule
module XOR3D1 (A1, A2, A3, Z);
  input A1, A2, A3;
  output Z;
endmodule
module XOR3D2 (A1, A2, A3, Z);
  input A1, A2, A3;
  output Z;
endmodule
module XOR3D4 (A1, A2, A3, Z);
  input A1, A2, A3;
  output Z;
endmodule
module XOR4D0 (A1, A2, A3, A4, Z);
  input 	A1, A2, A3, A4;
  output 	Z;
endmodule
module XOR4D1 (A1, A2, A3, A4, Z);
  input 	A1, A2, A3, A4;
  output 	Z;
endmodule
module XOR4D2 (A1, A2, A3, A4, Z);
  input 	A1, A2, A3, A4;
  output 	Z;
endmodule
module XOR4D4 (A1, A2, A3, A4, Z);
  input 	A1, A2, A3, A4;
  output 	Z;
endmodule
module ISOHID1 (ISO, I, Z);
    input ISO, I;
    output Z;
endmodule
module ISOHID2 (ISO, I, Z);
    input ISO, I;
    output Z;
endmodule
module ISOHID4 (ISO, I, Z);
    input ISO, I;
    output Z;
endmodule
module ISOHID8 (ISO, I, Z);
    input ISO, I;
    output Z;
endmodule
module ISOLOD1 (ISO, I, Z);
    input ISO, I;
    output Z;
endmodule
module ISOLOD2 (ISO, I, Z);
    input ISO, I;
    output Z;
endmodule
module ISOLOD4 (ISO, I, Z);
    input ISO, I;
    output Z;
endmodule
module ISOLOD8 (ISO, I, Z);
    input ISO, I;
    output Z;
endmodule
module LVLHLD1 (I, Z);
    input I;
    output Z;
endmodule
module LVLHLD2 (I, Z);
    input I;
    output Z;
endmodule
module LVLHLD4 (I, Z);
    input I;
    output Z;
endmodule
module LVLHLD8 (I, Z);
    input I;
    output Z;
endmodule
module LVLLHCD1 (I, NSLEEP, Z);
    input I, NSLEEP;
    output Z;
endmodule
module LVLLHCD2 (I, NSLEEP, Z);
    input I, NSLEEP;
    output Z;
endmodule
module LVLLHCD4 (I, NSLEEP, Z);
    input I, NSLEEP;
    output Z;
endmodule
module LVLLHCD8 (I, NSLEEP, Z);
    input I, NSLEEP;
    output Z;
endmodule
module LVLLHD1 (I, Z);
    input I;
    output Z;
endmodule
module LVLLHD2 (I, Z);
    input I;
    output Z;
endmodule
module LVLLHD4 (I, Z);
    input I;
    output Z;
endmodule
module LVLLHD8 (I, Z);
    input I;
    output Z;
endmodule
module LVLLHFACD1 (I, NSLEEP, Z);
    input I, NSLEEP;
    output Z;
endmodule
module LVLLHFACD2 (I, NSLEEP, Z);
    input I, NSLEEP;
    output Z;
endmodule
module LVLLHFACD4 (I, NSLEEP, Z);
    input I, NSLEEP;
    output Z;
endmodule
module LVLLHFACD8 (I, NSLEEP, Z);
    input I, NSLEEP;
    output Z;
endmodule
module LVLLHFAD1 (I, Z);
    input I;
    output Z;
endmodule
module LVLLHFAD2 (I, Z);
    input I;
    output Z;
endmodule
module LVLLHFAD4 (I, Z);
    input I;
    output Z;
endmodule
module LVLLHFAD8 (I, Z);
    input I;
    output Z;
endmodule

