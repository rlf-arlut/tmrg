`default_nettype none
`timescale 1ns / 1ps

module test(input wire i, output wire z);
  assign z=i;
endmodule
