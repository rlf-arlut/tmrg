module test;
  function automatic mux;
  endfunction
endmodule

